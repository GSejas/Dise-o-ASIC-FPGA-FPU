/******************************************************************************
 * File	Name			: ks233.v
 * Package Module Name	: Elliptic Curve Cryptoprocessor for GF(2^233)
 * Author		    	: Chester Rebeiro
 * Date of Creation		: 1/Apr/2008
 * Type	of file			: Verilog source code
 * Synopsis			    : Automatically generated code for karatsuba 233 bit
 ******************************************************************************/


`ifndef __KS_233_V__
`define __KS_233_V__
//`include "ks117.v"
//`include "ks116.v"
module ks233(a, b, d);

input wire [232:0] a;
input wire [232:0] b;
output wire [464:0] d;

wire [230:0] m1;
wire [232:0] m2;
wire [232:0] m3;
wire [116:0] ahl;
wire [116:0] bhl;

ks117 ksm1(a[116:0], b[116:0], m2);
ks116 ksm2(a[232:117], b[232:117], m1);
assign ahl[115:0] = a[232:117] ^ a[115:0];
assign ahl[116] = a[116];
assign bhl[115:0] = b[232:117] ^ b[115:0];
assign bhl[116] = b[116];
ks117 ksm3(ahl, bhl, m3);

assign  d[00] = m2[00];   
assign  d[01] = m2[01];   
assign  d[02] = m2[02];   
assign  d[03] = m2[03];   
assign  d[04] = m2[04];   
assign  d[05] = m2[05];   
assign  d[06] = m2[06];   
assign  d[07] = m2[07];   
assign  d[08] = m2[08];   
assign  d[09] = m2[09];   
assign  d[10] = m2[10];   
assign  d[11] = m2[11];   
assign  d[12] = m2[12];   
assign  d[13] = m2[13];   
assign  d[14] = m2[14];   
assign  d[15] = m2[15];   
assign  d[16] = m2[16];   
assign  d[17] = m2[17];   
assign  d[18] = m2[18];   
assign  d[19] = m2[19];   
assign  d[20] = m2[20];   
assign  d[21] = m2[21];   
assign  d[22] = m2[22];   
assign  d[23] = m2[23];   
assign  d[24] = m2[24];   
assign  d[25] = m2[25];   
assign  d[26] = m2[26];   
assign  d[27] = m2[27];   
assign  d[28] = m2[28];   
assign  d[29] = m2[29];   
assign  d[30] = m2[30];   
assign  d[31] = m2[31];   
assign  d[32] = m2[32];   
assign  d[33] = m2[33];   
assign  d[34] = m2[34];   
assign  d[35] = m2[35];   
assign  d[36] = m2[36];   
assign  d[37] = m2[37];   
assign  d[38] = m2[38];   
assign  d[39] = m2[39];   
assign  d[40] = m2[40];   
assign  d[41] = m2[41];   
assign  d[42] = m2[42];   
assign  d[43] = m2[43];   
assign  d[44] = m2[44];   
assign  d[45] = m2[45];   
assign  d[46] = m2[46];   
assign  d[47] = m2[47];   
assign  d[48] = m2[48];   
assign  d[49] = m2[49];   
assign  d[50] = m2[50];   
assign  d[51] = m2[51];   
assign  d[52] = m2[52];   
assign  d[53] = m2[53];   
assign  d[54] = m2[54];   
assign  d[55] = m2[55];   
assign  d[56] = m2[56];   
assign  d[57] = m2[57];   
assign  d[58] = m2[58];   
assign  d[59] = m2[59];   
assign  d[60] = m2[60];   
assign  d[61] = m2[61];   
assign  d[62] = m2[62];   
assign  d[63] = m2[63];   
assign  d[64] = m2[64];   
assign  d[65] = m2[65];   
assign  d[66] = m2[66];   
assign  d[67] = m2[67];   
assign  d[68] = m2[68];   
assign  d[69] = m2[69];   
assign  d[70] = m2[70];   
assign  d[71] = m2[71];   
assign  d[72] = m2[72];   
assign  d[73] = m2[73];   
assign  d[74] = m2[74];   
assign  d[75] = m2[75];   
assign  d[76] = m2[76];   
assign  d[77] = m2[77];   
assign  d[78] = m2[78];   
assign  d[79] = m2[79];   
assign  d[80] = m2[80];   
assign  d[81] = m2[81];   
assign  d[82] = m2[82];   
assign  d[83] = m2[83];   
assign  d[84] = m2[84];   
assign  d[85] = m2[85];   
assign  d[86] = m2[86];   
assign  d[87] = m2[87];   
assign  d[88] = m2[88];   
assign  d[89] = m2[89];   
assign  d[90] = m2[90];   
assign  d[91] = m2[91];   
assign  d[92] = m2[92];   
assign  d[93] = m2[93];   
assign  d[94] = m2[94];   
assign  d[95] = m2[95];   
assign  d[96] = m2[96];   
assign  d[97] = m2[97];   
assign  d[98] = m2[98];   
assign  d[99] = m2[99];   
assign  d[100] = m2[100];   
assign  d[101] = m2[101];   
assign  d[102] = m2[102];   
assign  d[103] = m2[103];   
assign  d[104] = m2[104];   
assign  d[105] = m2[105];   
assign  d[106] = m2[106];   
assign  d[107] = m2[107];   
assign  d[108] = m2[108];   
assign  d[109] = m2[109];   
assign  d[110] = m2[110];   
assign  d[111] = m2[111];   
assign  d[112] = m2[112];   
assign  d[113] = m2[113];   
assign  d[114] = m2[114];   
assign  d[115] = m2[115];   
assign  d[116] = m2[116];   
assign  d[117] = m2[117] ^ m1[00] ^ m2[00] ^ m3[00];   
assign  d[118] = m2[118] ^ m1[01] ^ m2[01] ^ m3[01];   
assign  d[119] = m2[119] ^ m1[02] ^ m2[02] ^ m3[02];   
assign  d[120] = m2[120] ^ m1[03] ^ m2[03] ^ m3[03];   
assign  d[121] = m2[121] ^ m1[04] ^ m2[04] ^ m3[04];   
assign  d[122] = m2[122] ^ m1[05] ^ m2[05] ^ m3[05];   
assign  d[123] = m2[123] ^ m1[06] ^ m2[06] ^ m3[06];   
assign  d[124] = m2[124] ^ m1[07] ^ m2[07] ^ m3[07];   
assign  d[125] = m2[125] ^ m1[08] ^ m2[08] ^ m3[08];   
assign  d[126] = m2[126] ^ m1[09] ^ m2[09] ^ m3[09];   
assign  d[127] = m2[127] ^ m1[10] ^ m2[10] ^ m3[10];   
assign  d[128] = m2[128] ^ m1[11] ^ m2[11] ^ m3[11];   
assign  d[129] = m2[129] ^ m1[12] ^ m2[12] ^ m3[12];   
assign  d[130] = m2[130] ^ m1[13] ^ m2[13] ^ m3[13];   
assign  d[131] = m2[131] ^ m1[14] ^ m2[14] ^ m3[14];   
assign  d[132] = m2[132] ^ m1[15] ^ m2[15] ^ m3[15];   
assign  d[133] = m2[133] ^ m1[16] ^ m2[16] ^ m3[16];   
assign  d[134] = m2[134] ^ m1[17] ^ m2[17] ^ m3[17];   
assign  d[135] = m2[135] ^ m1[18] ^ m2[18] ^ m3[18];   
assign  d[136] = m2[136] ^ m1[19] ^ m2[19] ^ m3[19];   
assign  d[137] = m2[137] ^ m1[20] ^ m2[20] ^ m3[20];   
assign  d[138] = m2[138] ^ m1[21] ^ m2[21] ^ m3[21];   
assign  d[139] = m2[139] ^ m1[22] ^ m2[22] ^ m3[22];   
assign  d[140] = m2[140] ^ m1[23] ^ m2[23] ^ m3[23];   
assign  d[141] = m2[141] ^ m1[24] ^ m2[24] ^ m3[24];   
assign  d[142] = m2[142] ^ m1[25] ^ m2[25] ^ m3[25];   
assign  d[143] = m2[143] ^ m1[26] ^ m2[26] ^ m3[26];   
assign  d[144] = m2[144] ^ m1[27] ^ m2[27] ^ m3[27];   
assign  d[145] = m2[145] ^ m1[28] ^ m2[28] ^ m3[28];   
assign  d[146] = m2[146] ^ m1[29] ^ m2[29] ^ m3[29];   
assign  d[147] = m2[147] ^ m1[30] ^ m2[30] ^ m3[30];   
assign  d[148] = m2[148] ^ m1[31] ^ m2[31] ^ m3[31];   
assign  d[149] = m2[149] ^ m1[32] ^ m2[32] ^ m3[32];   
assign  d[150] = m2[150] ^ m1[33] ^ m2[33] ^ m3[33];   
assign  d[151] = m2[151] ^ m1[34] ^ m2[34] ^ m3[34];   
assign  d[152] = m2[152] ^ m1[35] ^ m2[35] ^ m3[35];   
assign  d[153] = m2[153] ^ m1[36] ^ m2[36] ^ m3[36];   
assign  d[154] = m2[154] ^ m1[37] ^ m2[37] ^ m3[37];   
assign  d[155] = m2[155] ^ m1[38] ^ m2[38] ^ m3[38];   
assign  d[156] = m2[156] ^ m1[39] ^ m2[39] ^ m3[39];   
assign  d[157] = m2[157] ^ m1[40] ^ m2[40] ^ m3[40];   
assign  d[158] = m2[158] ^ m1[41] ^ m2[41] ^ m3[41];   
assign  d[159] = m2[159] ^ m1[42] ^ m2[42] ^ m3[42];   
assign  d[160] = m2[160] ^ m1[43] ^ m2[43] ^ m3[43];   
assign  d[161] = m2[161] ^ m1[44] ^ m2[44] ^ m3[44];   
assign  d[162] = m2[162] ^ m1[45] ^ m2[45] ^ m3[45];   
assign  d[163] = m2[163] ^ m1[46] ^ m2[46] ^ m3[46];   
assign  d[164] = m2[164] ^ m1[47] ^ m2[47] ^ m3[47];   
assign  d[165] = m2[165] ^ m1[48] ^ m2[48] ^ m3[48];   
assign  d[166] = m2[166] ^ m1[49] ^ m2[49] ^ m3[49];   
assign  d[167] = m2[167] ^ m1[50] ^ m2[50] ^ m3[50];   
assign  d[168] = m2[168] ^ m1[51] ^ m2[51] ^ m3[51];   
assign  d[169] = m2[169] ^ m1[52] ^ m2[52] ^ m3[52];   
assign  d[170] = m2[170] ^ m1[53] ^ m2[53] ^ m3[53];   
assign  d[171] = m2[171] ^ m1[54] ^ m2[54] ^ m3[54];   
assign  d[172] = m2[172] ^ m1[55] ^ m2[55] ^ m3[55];   
assign  d[173] = m2[173] ^ m1[56] ^ m2[56] ^ m3[56];   
assign  d[174] = m2[174] ^ m1[57] ^ m2[57] ^ m3[57];   
assign  d[175] = m2[175] ^ m1[58] ^ m2[58] ^ m3[58];   
assign  d[176] = m2[176] ^ m1[59] ^ m2[59] ^ m3[59];   
assign  d[177] = m2[177] ^ m1[60] ^ m2[60] ^ m3[60];   
assign  d[178] = m2[178] ^ m1[61] ^ m2[61] ^ m3[61];   
assign  d[179] = m2[179] ^ m1[62] ^ m2[62] ^ m3[62];   
assign  d[180] = m2[180] ^ m1[63] ^ m2[63] ^ m3[63];   
assign  d[181] = m2[181] ^ m1[64] ^ m2[64] ^ m3[64];   
assign  d[182] = m2[182] ^ m1[65] ^ m2[65] ^ m3[65];   
assign  d[183] = m2[183] ^ m1[66] ^ m2[66] ^ m3[66];   
assign  d[184] = m2[184] ^ m1[67] ^ m2[67] ^ m3[67];   
assign  d[185] = m2[185] ^ m1[68] ^ m2[68] ^ m3[68];   
assign  d[186] = m2[186] ^ m1[69] ^ m2[69] ^ m3[69];   
assign  d[187] = m2[187] ^ m1[70] ^ m2[70] ^ m3[70];   
assign  d[188] = m2[188] ^ m1[71] ^ m2[71] ^ m3[71];   
assign  d[189] = m2[189] ^ m1[72] ^ m2[72] ^ m3[72];   
assign  d[190] = m2[190] ^ m1[73] ^ m2[73] ^ m3[73];   
assign  d[191] = m2[191] ^ m1[74] ^ m2[74] ^ m3[74];   
assign  d[192] = m2[192] ^ m1[75] ^ m2[75] ^ m3[75];   
assign  d[193] = m2[193] ^ m1[76] ^ m2[76] ^ m3[76];   
assign  d[194] = m2[194] ^ m1[77] ^ m2[77] ^ m3[77];   
assign  d[195] = m2[195] ^ m1[78] ^ m2[78] ^ m3[78];   
assign  d[196] = m2[196] ^ m1[79] ^ m2[79] ^ m3[79];   
assign  d[197] = m2[197] ^ m1[80] ^ m2[80] ^ m3[80];   
assign  d[198] = m2[198] ^ m1[81] ^ m2[81] ^ m3[81];   
assign  d[199] = m2[199] ^ m1[82] ^ m2[82] ^ m3[82];   
assign  d[200] = m2[200] ^ m1[83] ^ m2[83] ^ m3[83];   
assign  d[201] = m2[201] ^ m1[84] ^ m2[84] ^ m3[84];   
assign  d[202] = m2[202] ^ m1[85] ^ m2[85] ^ m3[85];   
assign  d[203] = m2[203] ^ m1[86] ^ m2[86] ^ m3[86];   
assign  d[204] = m2[204] ^ m1[87] ^ m2[87] ^ m3[87];   
assign  d[205] = m2[205] ^ m1[88] ^ m2[88] ^ m3[88];   
assign  d[206] = m2[206] ^ m1[89] ^ m2[89] ^ m3[89];   
assign  d[207] = m2[207] ^ m1[90] ^ m2[90] ^ m3[90];   
assign  d[208] = m2[208] ^ m1[91] ^ m2[91] ^ m3[91];   
assign  d[209] = m2[209] ^ m1[92] ^ m2[92] ^ m3[92];   
assign  d[210] = m2[210] ^ m1[93] ^ m2[93] ^ m3[93];   
assign  d[211] = m2[211] ^ m1[94] ^ m2[94] ^ m3[94];   
assign  d[212] = m2[212] ^ m1[95] ^ m2[95] ^ m3[95];   
assign  d[213] = m2[213] ^ m1[96] ^ m2[96] ^ m3[96];   
assign  d[214] = m2[214] ^ m1[97] ^ m2[97] ^ m3[97];   
assign  d[215] = m2[215] ^ m1[98] ^ m2[98] ^ m3[98];   
assign  d[216] = m2[216] ^ m1[99] ^ m2[99] ^ m3[99];   
assign  d[217] = m2[217] ^ m1[100] ^ m2[100] ^ m3[100];   
assign  d[218] = m2[218] ^ m1[101] ^ m2[101] ^ m3[101];   
assign  d[219] = m2[219] ^ m1[102] ^ m2[102] ^ m3[102];   
assign  d[220] = m2[220] ^ m1[103] ^ m2[103] ^ m3[103];   
assign  d[221] = m2[221] ^ m1[104] ^ m2[104] ^ m3[104];   
assign  d[222] = m2[222] ^ m1[105] ^ m2[105] ^ m3[105];   
assign  d[223] = m2[223] ^ m1[106] ^ m2[106] ^ m3[106];   
assign  d[224] = m2[224] ^ m1[107] ^ m2[107] ^ m3[107];   
assign  d[225] = m2[225] ^ m1[108] ^ m2[108] ^ m3[108];   
assign  d[226] = m2[226] ^ m1[109] ^ m2[109] ^ m3[109];   
assign  d[227] = m2[227] ^ m1[110] ^ m2[110] ^ m3[110];   
assign  d[228] = m2[228] ^ m1[111] ^ m2[111] ^ m3[111];   
assign  d[229] = m2[229] ^ m1[112] ^ m2[112] ^ m3[112];   
assign  d[230] = m2[230] ^ m1[113] ^ m2[113] ^ m3[113];   
assign  d[231] = m2[231] ^ m1[114] ^ m2[114] ^ m3[114];   
assign  d[232] = m2[232] ^ m1[115] ^ m2[115] ^ m3[115];   
assign  d[233] = m1[116] ^ m2[116] ^ m3[116];   
assign  d[234] = m1[117] ^ m2[117] ^ m3[117] ^ m1[00];   
assign  d[235] = m1[118] ^ m2[118] ^ m3[118] ^ m1[01];   
assign  d[236] = m1[119] ^ m2[119] ^ m3[119] ^ m1[02];   
assign  d[237] = m1[120] ^ m2[120] ^ m3[120] ^ m1[03];   
assign  d[238] = m1[121] ^ m2[121] ^ m3[121] ^ m1[04];   
assign  d[239] = m1[122] ^ m2[122] ^ m3[122] ^ m1[05];   
assign  d[240] = m1[123] ^ m2[123] ^ m3[123] ^ m1[06];   
assign  d[241] = m1[124] ^ m2[124] ^ m3[124] ^ m1[07];   
assign  d[242] = m1[125] ^ m2[125] ^ m3[125] ^ m1[08];   
assign  d[243] = m1[126] ^ m2[126] ^ m3[126] ^ m1[09];   
assign  d[244] = m1[127] ^ m2[127] ^ m3[127] ^ m1[10];   
assign  d[245] = m1[128] ^ m2[128] ^ m3[128] ^ m1[11];   
assign  d[246] = m1[129] ^ m2[129] ^ m3[129] ^ m1[12];   
assign  d[247] = m1[130] ^ m2[130] ^ m3[130] ^ m1[13];   
assign  d[248] = m1[131] ^ m2[131] ^ m3[131] ^ m1[14];   
assign  d[249] = m1[132] ^ m2[132] ^ m3[132] ^ m1[15];   
assign  d[250] = m1[133] ^ m2[133] ^ m3[133] ^ m1[16];   
assign  d[251] = m1[134] ^ m2[134] ^ m3[134] ^ m1[17];   
assign  d[252] = m1[135] ^ m2[135] ^ m3[135] ^ m1[18];   
assign  d[253] = m1[136] ^ m2[136] ^ m3[136] ^ m1[19];   
assign  d[254] = m1[137] ^ m2[137] ^ m3[137] ^ m1[20];   
assign  d[255] = m1[138] ^ m2[138] ^ m3[138] ^ m1[21];   
assign  d[256] = m1[139] ^ m2[139] ^ m3[139] ^ m1[22];   
assign  d[257] = m1[140] ^ m2[140] ^ m3[140] ^ m1[23];   
assign  d[258] = m1[141] ^ m2[141] ^ m3[141] ^ m1[24];   
assign  d[259] = m1[142] ^ m2[142] ^ m3[142] ^ m1[25];   
assign  d[260] = m1[143] ^ m2[143] ^ m3[143] ^ m1[26];   
assign  d[261] = m1[144] ^ m2[144] ^ m3[144] ^ m1[27];   
assign  d[262] = m1[145] ^ m2[145] ^ m3[145] ^ m1[28];   
assign  d[263] = m1[146] ^ m2[146] ^ m3[146] ^ m1[29];   
assign  d[264] = m1[147] ^ m2[147] ^ m3[147] ^ m1[30];   
assign  d[265] = m1[148] ^ m2[148] ^ m3[148] ^ m1[31];   
assign  d[266] = m1[149] ^ m2[149] ^ m3[149] ^ m1[32];   
assign  d[267] = m1[150] ^ m2[150] ^ m3[150] ^ m1[33];   
assign  d[268] = m1[151] ^ m2[151] ^ m3[151] ^ m1[34];   
assign  d[269] = m1[152] ^ m2[152] ^ m3[152] ^ m1[35];   
assign  d[270] = m1[153] ^ m2[153] ^ m3[153] ^ m1[36];   
assign  d[271] = m1[154] ^ m2[154] ^ m3[154] ^ m1[37];   
assign  d[272] = m1[155] ^ m2[155] ^ m3[155] ^ m1[38];   
assign  d[273] = m1[156] ^ m2[156] ^ m3[156] ^ m1[39];   
assign  d[274] = m1[157] ^ m2[157] ^ m3[157] ^ m1[40];   
assign  d[275] = m1[158] ^ m2[158] ^ m3[158] ^ m1[41];   
assign  d[276] = m1[159] ^ m2[159] ^ m3[159] ^ m1[42];   
assign  d[277] = m1[160] ^ m2[160] ^ m3[160] ^ m1[43];   
assign  d[278] = m1[161] ^ m2[161] ^ m3[161] ^ m1[44];   
assign  d[279] = m1[162] ^ m2[162] ^ m3[162] ^ m1[45];   
assign  d[280] = m1[163] ^ m2[163] ^ m3[163] ^ m1[46];   
assign  d[281] = m1[164] ^ m2[164] ^ m3[164] ^ m1[47];   
assign  d[282] = m1[165] ^ m2[165] ^ m3[165] ^ m1[48];   
assign  d[283] = m1[166] ^ m2[166] ^ m3[166] ^ m1[49];   
assign  d[284] = m1[167] ^ m2[167] ^ m3[167] ^ m1[50];   
assign  d[285] = m1[168] ^ m2[168] ^ m3[168] ^ m1[51];   
assign  d[286] = m1[169] ^ m2[169] ^ m3[169] ^ m1[52];   
assign  d[287] = m1[170] ^ m2[170] ^ m3[170] ^ m1[53];   
assign  d[288] = m1[171] ^ m2[171] ^ m3[171] ^ m1[54];   
assign  d[289] = m1[172] ^ m2[172] ^ m3[172] ^ m1[55];   
assign  d[290] = m1[173] ^ m2[173] ^ m3[173] ^ m1[56];   
assign  d[291] = m1[174] ^ m2[174] ^ m3[174] ^ m1[57];   
assign  d[292] = m1[175] ^ m2[175] ^ m3[175] ^ m1[58];   
assign  d[293] = m1[176] ^ m2[176] ^ m3[176] ^ m1[59];   
assign  d[294] = m1[177] ^ m2[177] ^ m3[177] ^ m1[60];   
assign  d[295] = m1[178] ^ m2[178] ^ m3[178] ^ m1[61];   
assign  d[296] = m1[179] ^ m2[179] ^ m3[179] ^ m1[62];   
assign  d[297] = m1[180] ^ m2[180] ^ m3[180] ^ m1[63];   
assign  d[298] = m1[181] ^ m2[181] ^ m3[181] ^ m1[64];   
assign  d[299] = m1[182] ^ m2[182] ^ m3[182] ^ m1[65];   
assign  d[300] = m1[183] ^ m2[183] ^ m3[183] ^ m1[66];   
assign  d[301] = m1[184] ^ m2[184] ^ m3[184] ^ m1[67];   
assign  d[302] = m1[185] ^ m2[185] ^ m3[185] ^ m1[68];   
assign  d[303] = m1[186] ^ m2[186] ^ m3[186] ^ m1[69];   
assign  d[304] = m1[187] ^ m2[187] ^ m3[187] ^ m1[70];   
assign  d[305] = m1[188] ^ m2[188] ^ m3[188] ^ m1[71];   
assign  d[306] = m1[189] ^ m2[189] ^ m3[189] ^ m1[72];   
assign  d[307] = m1[190] ^ m2[190] ^ m3[190] ^ m1[73];   
assign  d[308] = m1[191] ^ m2[191] ^ m3[191] ^ m1[74];   
assign  d[309] = m1[192] ^ m2[192] ^ m3[192] ^ m1[75];   
assign  d[310] = m1[193] ^ m2[193] ^ m3[193] ^ m1[76];   
assign  d[311] = m1[194] ^ m2[194] ^ m3[194] ^ m1[77];   
assign  d[312] = m1[195] ^ m2[195] ^ m3[195] ^ m1[78];   
assign  d[313] = m1[196] ^ m2[196] ^ m3[196] ^ m1[79];   
assign  d[314] = m1[197] ^ m2[197] ^ m3[197] ^ m1[80];   
assign  d[315] = m1[198] ^ m2[198] ^ m3[198] ^ m1[81];   
assign  d[316] = m1[199] ^ m2[199] ^ m3[199] ^ m1[82];   
assign  d[317] = m1[200] ^ m2[200] ^ m3[200] ^ m1[83];   
assign  d[318] = m1[201] ^ m2[201] ^ m3[201] ^ m1[84];   
assign  d[319] = m1[202] ^ m2[202] ^ m3[202] ^ m1[85];   
assign  d[320] = m1[203] ^ m2[203] ^ m3[203] ^ m1[86];   
assign  d[321] = m1[204] ^ m2[204] ^ m3[204] ^ m1[87];   
assign  d[322] = m1[205] ^ m2[205] ^ m3[205] ^ m1[88];   
assign  d[323] = m1[206] ^ m2[206] ^ m3[206] ^ m1[89];   
assign  d[324] = m1[207] ^ m2[207] ^ m3[207] ^ m1[90];   
assign  d[325] = m1[208] ^ m2[208] ^ m3[208] ^ m1[91];   
assign  d[326] = m1[209] ^ m2[209] ^ m3[209] ^ m1[92];   
assign  d[327] = m1[210] ^ m2[210] ^ m3[210] ^ m1[93];   
assign  d[328] = m1[211] ^ m2[211] ^ m3[211] ^ m1[94];   
assign  d[329] = m1[212] ^ m2[212] ^ m3[212] ^ m1[95];   
assign  d[330] = m1[213] ^ m2[213] ^ m3[213] ^ m1[96];   
assign  d[331] = m1[214] ^ m2[214] ^ m3[214] ^ m1[97];   
assign  d[332] = m1[215] ^ m2[215] ^ m3[215] ^ m1[98];   
assign  d[333] = m1[216] ^ m2[216] ^ m3[216] ^ m1[99];   
assign  d[334] = m1[217] ^ m2[217] ^ m3[217] ^ m1[100];   
assign  d[335] = m1[218] ^ m2[218] ^ m3[218] ^ m1[101];   
assign  d[336] = m1[219] ^ m2[219] ^ m3[219] ^ m1[102];   
assign  d[337] = m1[220] ^ m2[220] ^ m3[220] ^ m1[103];   
assign  d[338] = m1[221] ^ m2[221] ^ m3[221] ^ m1[104];   
assign  d[339] = m1[222] ^ m2[222] ^ m3[222] ^ m1[105];   
assign  d[340] = m1[223] ^ m2[223] ^ m3[223] ^ m1[106];   
assign  d[341] = m1[224] ^ m2[224] ^ m3[224] ^ m1[107];   
assign  d[342] = m1[225] ^ m2[225] ^ m3[225] ^ m1[108];   
assign  d[343] = m1[226] ^ m2[226] ^ m3[226] ^ m1[109];   
assign  d[344] = m1[227] ^ m2[227] ^ m3[227] ^ m1[110];   
assign  d[345] = m1[228] ^ m2[228] ^ m3[228] ^ m1[111];   
assign  d[346] = m1[229] ^ m2[229] ^ m3[229] ^ m1[112];   
assign  d[347] = m1[230] ^ m2[230] ^ m3[230] ^ m1[113];   
assign  d[348] = m2[231] ^ m3[231] ^ m1[114];   
assign  d[349] = m2[232] ^ m3[232] ^ m1[115];   
assign  d[350] = m1[116];   
assign  d[351] = m1[117];   
assign  d[352] = m1[118];   
assign  d[353] = m1[119];   
assign  d[354] = m1[120];   
assign  d[355] = m1[121];   
assign  d[356] = m1[122];   
assign  d[357] = m1[123];   
assign  d[358] = m1[124];   
assign  d[359] = m1[125];   
assign  d[360] = m1[126];   
assign  d[361] = m1[127];   
assign  d[362] = m1[128];   
assign  d[363] = m1[129];   
assign  d[364] = m1[130];   
assign  d[365] = m1[131];   
assign  d[366] = m1[132];   
assign  d[367] = m1[133];   
assign  d[368] = m1[134];   
assign  d[369] = m1[135];   
assign  d[370] = m1[136];   
assign  d[371] = m1[137];   
assign  d[372] = m1[138];   
assign  d[373] = m1[139];   
assign  d[374] = m1[140];   
assign  d[375] = m1[141];   
assign  d[376] = m1[142];   
assign  d[377] = m1[143];   
assign  d[378] = m1[144];   
assign  d[379] = m1[145];   
assign  d[380] = m1[146];   
assign  d[381] = m1[147];   
assign  d[382] = m1[148];   
assign  d[383] = m1[149];   
assign  d[384] = m1[150];   
assign  d[385] = m1[151];   
assign  d[386] = m1[152];   
assign  d[387] = m1[153];   
assign  d[388] = m1[154];   
assign  d[389] = m1[155];   
assign  d[390] = m1[156];   
assign  d[391] = m1[157];   
assign  d[392] = m1[158];   
assign  d[393] = m1[159];   
assign  d[394] = m1[160];   
assign  d[395] = m1[161];   
assign  d[396] = m1[162];   
assign  d[397] = m1[163];   
assign  d[398] = m1[164];   
assign  d[399] = m1[165];   
assign  d[400] = m1[166];   
assign  d[401] = m1[167];   
assign  d[402] = m1[168];   
assign  d[403] = m1[169];   
assign  d[404] = m1[170];   
assign  d[405] = m1[171];   
assign  d[406] = m1[172];   
assign  d[407] = m1[173];   
assign  d[408] = m1[174];   
assign  d[409] = m1[175];   
assign  d[410] = m1[176];   
assign  d[411] = m1[177];   
assign  d[412] = m1[178];   
assign  d[413] = m1[179];   
assign  d[414] = m1[180];   
assign  d[415] = m1[181];   
assign  d[416] = m1[182];   
assign  d[417] = m1[183];   
assign  d[418] = m1[184];   
assign  d[419] = m1[185];   
assign  d[420] = m1[186];   
assign  d[421] = m1[187];   
assign  d[422] = m1[188];   
assign  d[423] = m1[189];   
assign  d[424] = m1[190];   
assign  d[425] = m1[191];   
assign  d[426] = m1[192];   
assign  d[427] = m1[193];   
assign  d[428] = m1[194];   
assign  d[429] = m1[195];   
assign  d[430] = m1[196];   
assign  d[431] = m1[197];   
assign  d[432] = m1[198];   
assign  d[433] = m1[199];   
assign  d[434] = m1[200];   
assign  d[435] = m1[201];   
assign  d[436] = m1[202];   
assign  d[437] = m1[203];   
assign  d[438] = m1[204];   
assign  d[439] = m1[205];   
assign  d[440] = m1[206];   
assign  d[441] = m1[207];   
assign  d[442] = m1[208];   
assign  d[443] = m1[209];   
assign  d[444] = m1[210];   
assign  d[445] = m1[211];   
assign  d[446] = m1[212];   
assign  d[447] = m1[213];   
assign  d[448] = m1[214];   
assign  d[449] = m1[215];   
assign  d[450] = m1[216];   
assign  d[451] = m1[217];   
assign  d[452] = m1[218];   
assign  d[453] = m1[219];   
assign  d[454] = m1[220];   
assign  d[455] = m1[221];   
assign  d[456] = m1[222];   
assign  d[457] = m1[223];   
assign  d[458] = m1[224];   
assign  d[459] = m1[225];   
assign  d[460] = m1[226];   
assign  d[461] = m1[227];   
assign  d[462] = m1[228];   
assign  d[463] = m1[229];   
assign  d[464] = m1[230];   
endmodule
`endif
