/******************************************************************************
 * File	Name			: mod.v
 * Package Module Name	: Elliptic Curve Cryptoprocessor for GF(2^233)
 * Author		    	: Chester Rebeiro
 * Date of Creation		: 1/Apr/2008
 * Type	of file			: Verilog source code
 * Synopsis			    : Automatically generated code for modulo operation
 *  with the irreducible polynomial x^233 + x^74 + 1
 ******************************************************************************/

`ifndef __MOD_V__
`define __MOD_V__
module mod(a, d);

input wire [464:0] a;
output wire [232:0] d;

assign d[0] = a[0] ^ a[233] ^ a[392];
assign d[1] = a[1] ^ a[234] ^ a[393];
assign d[2] = a[2] ^ a[235] ^ a[394];
assign d[3] = a[3] ^ a[236] ^ a[395];
assign d[4] = a[4] ^ a[237] ^ a[396];
assign d[5] = a[5] ^ a[238] ^ a[397];
assign d[6] = a[6] ^ a[239] ^ a[398];
assign d[7] = a[7] ^ a[240] ^ a[399];
assign d[8] = a[8] ^ a[241] ^ a[400];
assign d[9] = a[9] ^ a[242] ^ a[401];
assign d[10] = a[10] ^ a[243] ^ a[402];
assign d[11] = a[11] ^ a[244] ^ a[403];
assign d[12] = a[12] ^ a[245] ^ a[404];
assign d[13] = a[13] ^ a[246] ^ a[405];
assign d[14] = a[14] ^ a[247] ^ a[406];
assign d[15] = a[15] ^ a[248] ^ a[407];
assign d[16] = a[16] ^ a[249] ^ a[408];
assign d[17] = a[17] ^ a[250] ^ a[409];
assign d[18] = a[18] ^ a[251] ^ a[410];
assign d[19] = a[19] ^ a[252] ^ a[411];
assign d[20] = a[20] ^ a[253] ^ a[412];
assign d[21] = a[21] ^ a[254] ^ a[413];
assign d[22] = a[22] ^ a[255] ^ a[414];
assign d[23] = a[23] ^ a[256] ^ a[415];
assign d[24] = a[24] ^ a[257] ^ a[416];
assign d[25] = a[25] ^ a[258] ^ a[417];
assign d[26] = a[26] ^ a[259] ^ a[418];
assign d[27] = a[27] ^ a[260] ^ a[419];
assign d[28] = a[28] ^ a[261] ^ a[420];
assign d[29] = a[29] ^ a[262] ^ a[421];
assign d[30] = a[30] ^ a[263] ^ a[422];
assign d[31] = a[31] ^ a[264] ^ a[423];
assign d[32] = a[32] ^ a[265] ^ a[424];
assign d[33] = a[33] ^ a[266] ^ a[425];
assign d[34] = a[34] ^ a[267] ^ a[426];
assign d[35] = a[35] ^ a[268] ^ a[427];
assign d[36] = a[36] ^ a[269] ^ a[428];
assign d[37] = a[37] ^ a[270] ^ a[429];
assign d[38] = a[38] ^ a[271] ^ a[430];
assign d[39] = a[39] ^ a[272] ^ a[431];
assign d[40] = a[40] ^ a[273] ^ a[432];
assign d[41] = a[41] ^ a[274] ^ a[433];
assign d[42] = a[42] ^ a[275] ^ a[434];
assign d[43] = a[43] ^ a[276] ^ a[435];
assign d[44] = a[44] ^ a[277] ^ a[436];
assign d[45] = a[45] ^ a[278] ^ a[437];
assign d[46] = a[46] ^ a[279] ^ a[438];
assign d[47] = a[47] ^ a[280] ^ a[439];
assign d[48] = a[48] ^ a[281] ^ a[440];
assign d[49] = a[49] ^ a[282] ^ a[441];
assign d[50] = a[50] ^ a[283] ^ a[442];
assign d[51] = a[51] ^ a[284] ^ a[443];
assign d[52] = a[52] ^ a[285] ^ a[444];
assign d[53] = a[53] ^ a[286] ^ a[445];
assign d[54] = a[54] ^ a[287] ^ a[446];
assign d[55] = a[55] ^ a[288] ^ a[447];
assign d[56] = a[56] ^ a[289] ^ a[448];
assign d[57] = a[57] ^ a[290] ^ a[449];
assign d[58] = a[58] ^ a[291] ^ a[450];
assign d[59] = a[59] ^ a[292] ^ a[451];
assign d[60] = a[60] ^ a[293] ^ a[452];
assign d[61] = a[61] ^ a[294] ^ a[453];
assign d[62] = a[62] ^ a[295] ^ a[454];
assign d[63] = a[63] ^ a[296] ^ a[455];
assign d[64] = a[64] ^ a[297] ^ a[456];
assign d[65] = a[65] ^ a[298] ^ a[457];
assign d[66] = a[66] ^ a[299] ^ a[458];
assign d[67] = a[67] ^ a[300] ^ a[459];
assign d[68] = a[68] ^ a[301] ^ a[460];
assign d[69] = a[69] ^ a[302] ^ a[461];
assign d[70] = a[70] ^ a[303] ^ a[462];
assign d[71] = a[71] ^ a[304] ^ a[463];
assign d[72] = a[72] ^ a[305] ^ a[464];
assign d[73] = a[73] ^ a[306];
assign d[74] = a[74] ^ a[233] ^ a[307] ^ a[392];
assign d[75] = a[75] ^ a[234] ^ a[308] ^ a[393];
assign d[76] = a[76] ^ a[235] ^ a[309] ^ a[394];
assign d[77] = a[77] ^ a[236] ^ a[310] ^ a[395];
assign d[78] = a[78] ^ a[237] ^ a[311] ^ a[396];
assign d[79] = a[79] ^ a[238] ^ a[312] ^ a[397];
assign d[80] = a[80] ^ a[239] ^ a[313] ^ a[398];
assign d[81] = a[81] ^ a[240] ^ a[314] ^ a[399];
assign d[82] = a[82] ^ a[241] ^ a[315] ^ a[400];
assign d[83] = a[83] ^ a[242] ^ a[316] ^ a[401];
assign d[84] = a[84] ^ a[243] ^ a[317] ^ a[402];
assign d[85] = a[85] ^ a[244] ^ a[318] ^ a[403];
assign d[86] = a[86] ^ a[245] ^ a[319] ^ a[404];
assign d[87] = a[87] ^ a[246] ^ a[320] ^ a[405];
assign d[88] = a[88] ^ a[247] ^ a[321] ^ a[406];
assign d[89] = a[89] ^ a[248] ^ a[322] ^ a[407];
assign d[90] = a[90] ^ a[249] ^ a[323] ^ a[408];
assign d[91] = a[91] ^ a[250] ^ a[324] ^ a[409];
assign d[92] = a[92] ^ a[251] ^ a[325] ^ a[410];
assign d[93] = a[93] ^ a[252] ^ a[326] ^ a[411];
assign d[94] = a[94] ^ a[253] ^ a[327] ^ a[412];
assign d[95] = a[95] ^ a[254] ^ a[328] ^ a[413];
assign d[96] = a[96] ^ a[255] ^ a[329] ^ a[414];
assign d[97] = a[97] ^ a[256] ^ a[330] ^ a[415];
assign d[98] = a[98] ^ a[257] ^ a[331] ^ a[416];
assign d[99] = a[99] ^ a[258] ^ a[332] ^ a[417];
assign d[100] = a[100] ^ a[259] ^ a[333] ^ a[418];
assign d[101] = a[101] ^ a[260] ^ a[334] ^ a[419];
assign d[102] = a[102] ^ a[261] ^ a[335] ^ a[420];
assign d[103] = a[103] ^ a[262] ^ a[336] ^ a[421];
assign d[104] = a[104] ^ a[263] ^ a[337] ^ a[422];
assign d[105] = a[105] ^ a[264] ^ a[338] ^ a[423];
assign d[106] = a[106] ^ a[265] ^ a[339] ^ a[424];
assign d[107] = a[107] ^ a[266] ^ a[340] ^ a[425];
assign d[108] = a[108] ^ a[267] ^ a[341] ^ a[426];
assign d[109] = a[109] ^ a[268] ^ a[342] ^ a[427];
assign d[110] = a[110] ^ a[269] ^ a[343] ^ a[428];
assign d[111] = a[111] ^ a[270] ^ a[344] ^ a[429];
assign d[112] = a[112] ^ a[271] ^ a[345] ^ a[430];
assign d[113] = a[113] ^ a[272] ^ a[346] ^ a[431];
assign d[114] = a[114] ^ a[273] ^ a[347] ^ a[432];
assign d[115] = a[115] ^ a[274] ^ a[348] ^ a[433];
assign d[116] = a[116] ^ a[275] ^ a[349] ^ a[434];
assign d[117] = a[117] ^ a[276] ^ a[350] ^ a[435];
assign d[118] = a[118] ^ a[277] ^ a[351] ^ a[436];
assign d[119] = a[119] ^ a[278] ^ a[352] ^ a[437];
assign d[120] = a[120] ^ a[279] ^ a[353] ^ a[438];
assign d[121] = a[121] ^ a[280] ^ a[354] ^ a[439];
assign d[122] = a[122] ^ a[281] ^ a[355] ^ a[440];
assign d[123] = a[123] ^ a[282] ^ a[356] ^ a[441];
assign d[124] = a[124] ^ a[283] ^ a[357] ^ a[442];
assign d[125] = a[125] ^ a[284] ^ a[358] ^ a[443];
assign d[126] = a[126] ^ a[285] ^ a[359] ^ a[444];
assign d[127] = a[127] ^ a[286] ^ a[360] ^ a[445];
assign d[128] = a[128] ^ a[287] ^ a[361] ^ a[446];
assign d[129] = a[129] ^ a[288] ^ a[362] ^ a[447];
assign d[130] = a[130] ^ a[289] ^ a[363] ^ a[448];
assign d[131] = a[131] ^ a[290] ^ a[364] ^ a[449];
assign d[132] = a[132] ^ a[291] ^ a[365] ^ a[450];
assign d[133] = a[133] ^ a[292] ^ a[366] ^ a[451];
assign d[134] = a[134] ^ a[293] ^ a[367] ^ a[452];
assign d[135] = a[135] ^ a[294] ^ a[368] ^ a[453];
assign d[136] = a[136] ^ a[295] ^ a[369] ^ a[454];
assign d[137] = a[137] ^ a[296] ^ a[370] ^ a[455];
assign d[138] = a[138] ^ a[297] ^ a[371] ^ a[456];
assign d[139] = a[139] ^ a[298] ^ a[372] ^ a[457];
assign d[140] = a[140] ^ a[299] ^ a[373] ^ a[458];
assign d[141] = a[141] ^ a[300] ^ a[374] ^ a[459];
assign d[142] = a[142] ^ a[301] ^ a[375] ^ a[460];
assign d[143] = a[143] ^ a[302] ^ a[376] ^ a[461];
assign d[144] = a[144] ^ a[303] ^ a[377] ^ a[462];
assign d[145] = a[145] ^ a[304] ^ a[378] ^ a[463];
assign d[146] = a[146] ^ a[305] ^ a[379] ^ a[464];
assign d[147] = a[147] ^ a[306] ^ a[380];
assign d[148] = a[148] ^ a[307] ^ a[381];
assign d[149] = a[149] ^ a[308] ^ a[382];
assign d[150] = a[150] ^ a[309] ^ a[383];
assign d[151] = a[151] ^ a[310] ^ a[384];
assign d[152] = a[152] ^ a[311] ^ a[385];
assign d[153] = a[153] ^ a[312] ^ a[386];
assign d[154] = a[154] ^ a[313] ^ a[387];
assign d[155] = a[155] ^ a[314] ^ a[388];
assign d[156] = a[156] ^ a[315] ^ a[389];
assign d[157] = a[157] ^ a[316] ^ a[390];
assign d[158] = a[158] ^ a[317] ^ a[391];
assign d[159] = a[159] ^ a[318] ^ a[392];
assign d[160] = a[160] ^ a[319] ^ a[393];
assign d[161] = a[161] ^ a[320] ^ a[394];
assign d[162] = a[162] ^ a[321] ^ a[395];
assign d[163] = a[163] ^ a[322] ^ a[396];
assign d[164] = a[164] ^ a[323] ^ a[397];
assign d[165] = a[165] ^ a[324] ^ a[398];
assign d[166] = a[166] ^ a[325] ^ a[399];
assign d[167] = a[167] ^ a[326] ^ a[400];
assign d[168] = a[168] ^ a[327] ^ a[401];
assign d[169] = a[169] ^ a[328] ^ a[402];
assign d[170] = a[170] ^ a[329] ^ a[403];
assign d[171] = a[171] ^ a[330] ^ a[404];
assign d[172] = a[172] ^ a[331] ^ a[405];
assign d[173] = a[173] ^ a[332] ^ a[406];
assign d[174] = a[174] ^ a[333] ^ a[407];
assign d[175] = a[175] ^ a[334] ^ a[408];
assign d[176] = a[176] ^ a[335] ^ a[409];
assign d[177] = a[177] ^ a[336] ^ a[410];
assign d[178] = a[178] ^ a[337] ^ a[411];
assign d[179] = a[179] ^ a[338] ^ a[412];
assign d[180] = a[180] ^ a[339] ^ a[413];
assign d[181] = a[181] ^ a[340] ^ a[414];
assign d[182] = a[182] ^ a[341] ^ a[415];
assign d[183] = a[183] ^ a[342] ^ a[416];
assign d[184] = a[184] ^ a[343] ^ a[417];
assign d[185] = a[185] ^ a[344] ^ a[418];
assign d[186] = a[186] ^ a[345] ^ a[419];
assign d[187] = a[187] ^ a[346] ^ a[420];
assign d[188] = a[188] ^ a[347] ^ a[421];
assign d[189] = a[189] ^ a[348] ^ a[422];
assign d[190] = a[190] ^ a[349] ^ a[423];
assign d[191] = a[191] ^ a[350] ^ a[424];
assign d[192] = a[192] ^ a[351] ^ a[425];
assign d[193] = a[193] ^ a[352] ^ a[426];
assign d[194] = a[194] ^ a[353] ^ a[427];
assign d[195] = a[195] ^ a[354] ^ a[428];
assign d[196] = a[196] ^ a[355] ^ a[429];
assign d[197] = a[197] ^ a[356] ^ a[430];
assign d[198] = a[198] ^ a[357] ^ a[431];
assign d[199] = a[199] ^ a[358] ^ a[432];
assign d[200] = a[200] ^ a[359] ^ a[433];
assign d[201] = a[201] ^ a[360] ^ a[434];
assign d[202] = a[202] ^ a[361] ^ a[435];
assign d[203] = a[203] ^ a[362] ^ a[436];
assign d[204] = a[204] ^ a[363] ^ a[437];
assign d[205] = a[205] ^ a[364] ^ a[438];
assign d[206] = a[206] ^ a[365] ^ a[439];
assign d[207] = a[207] ^ a[366] ^ a[440];
assign d[208] = a[208] ^ a[367] ^ a[441];
assign d[209] = a[209] ^ a[368] ^ a[442];
assign d[210] = a[210] ^ a[369] ^ a[443];
assign d[211] = a[211] ^ a[370] ^ a[444];
assign d[212] = a[212] ^ a[371] ^ a[445];
assign d[213] = a[213] ^ a[372] ^ a[446];
assign d[214] = a[214] ^ a[373] ^ a[447];
assign d[215] = a[215] ^ a[374] ^ a[448];
assign d[216] = a[216] ^ a[375] ^ a[449];
assign d[217] = a[217] ^ a[376] ^ a[450];
assign d[218] = a[218] ^ a[377] ^ a[451];
assign d[219] = a[219] ^ a[378] ^ a[452];
assign d[220] = a[220] ^ a[379] ^ a[453];
assign d[221] = a[221] ^ a[380] ^ a[454];
assign d[222] = a[222] ^ a[381] ^ a[455];
assign d[223] = a[223] ^ a[382] ^ a[456];
assign d[224] = a[224] ^ a[383] ^ a[457];
assign d[225] = a[225] ^ a[384] ^ a[458];
assign d[226] = a[226] ^ a[385] ^ a[459];
assign d[227] = a[227] ^ a[386] ^ a[460];
assign d[228] = a[228] ^ a[387] ^ a[461];
assign d[229] = a[229] ^ a[388] ^ a[462];
assign d[230] = a[230] ^ a[389] ^ a[463];
assign d[231] = a[231] ^ a[390] ^ a[464];
assign d[232] = a[232] ^ a[391];
endmodule
`endif
