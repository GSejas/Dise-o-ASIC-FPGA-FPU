LIBRARY ieee;
use IEEE.std_logic_1164.all;

package mdctrom2048 is

--n = 2048
constant rom_lenght_br: integer:=512;
constant rom_lenght: integer:=2560;
type rom_table is array (0 to rom_lenght-1) of std_logic_vector (31 downto 0);
type rom_bitrev is array (0 to rom_lenght_br-1) of std_logic_vector (31 downto 0);

constant bitrev: rom_bitrev:= rom_bitrev'(

X"000003fe",
X"00000000",
X"000001fe",
X"00000200",
X"000002fe",
X"00000100",
X"000000fe",
X"00000300",
X"0000037e",
X"00000080",
X"0000017e",
X"00000280",
X"0000027e",
X"00000180",
X"0000007e",
X"00000380",
X"000003be",
X"00000040",
X"000001be",
X"00000240",
X"000002be",
X"00000140",
X"000000be",
X"00000340",
X"0000033e",
X"000000c0",
X"0000013e",
X"000002c0",
X"0000023e",
X"000001c0",
X"0000003e",
X"000003c0",
X"000003de",
X"00000020",
X"000001de",
X"00000220",
X"000002de",
X"00000120",
X"000000de",
X"00000320",
X"0000035e",
X"000000a0",
X"0000015e",
X"000002a0",
X"0000025e",
X"000001a0",
X"0000005e",
X"000003a0",
X"0000039e",
X"00000060",
X"0000019e",
X"00000260",
X"0000029e",
X"00000160",
X"0000009e",
X"00000360",
X"0000031e",
X"000000e0",
X"0000011e",
X"000002e0",
X"0000021e",
X"000001e0",
X"0000001e",
X"000003e0",
X"000003ee",
X"00000010",
X"000001ee",
X"00000210",
X"000002ee",
X"00000110",
X"000000ee",
X"00000310",
X"0000036e",
X"00000090",
X"0000016e",
X"00000290",
X"0000026e",
X"00000190",
X"0000006e",
X"00000390",
X"000003ae",
X"00000050",
X"000001ae",
X"00000250",
X"000002ae",
X"00000150",
X"000000ae",
X"00000350",
X"0000032e",
X"000000d0",
X"0000012e",
X"000002d0",
X"0000022e",
X"000001d0",
X"0000002e",
X"000003d0",
X"000003ce",
X"00000030",
X"000001ce",
X"00000230",
X"000002ce",
X"00000130",
X"000000ce",
X"00000330",
X"0000034e",
X"000000b0",
X"0000014e",
X"000002b0",
X"0000024e",
X"000001b0",
X"0000004e",
X"000003b0",
X"0000038e",
X"00000070",
X"0000018e",
X"00000270",
X"0000028e",
X"00000170",
X"0000008e",
X"00000370",
X"0000030e",
X"000000f0",
X"0000010e",
X"000002f0",
X"0000020e",
X"000001f0",
X"0000000e",
X"000003f0",
X"000003f6",
X"00000008",
X"000001f6",
X"00000208",
X"000002f6",
X"00000108",
X"000000f6",
X"00000308",
X"00000376",
X"00000088",
X"00000176",
X"00000288",
X"00000276",
X"00000188",
X"00000076",
X"00000388",
X"000003b6",
X"00000048",
X"000001b6",
X"00000248",
X"000002b6",
X"00000148",
X"000000b6",
X"00000348",
X"00000336",
X"000000c8",
X"00000136",
X"000002c8",
X"00000236",
X"000001c8",
X"00000036",
X"000003c8",
X"000003d6",
X"00000028",
X"000001d6",
X"00000228",
X"000002d6",
X"00000128",
X"000000d6",
X"00000328",
X"00000356",
X"000000a8",
X"00000156",
X"000002a8",
X"00000256",
X"000001a8",
X"00000056",
X"000003a8",
X"00000396",
X"00000068",
X"00000196",
X"00000268",
X"00000296",
X"00000168",
X"00000096",
X"00000368",
X"00000316",
X"000000e8",
X"00000116",
X"000002e8",
X"00000216",
X"000001e8",
X"00000016",
X"000003e8",
X"000003e6",
X"00000018",
X"000001e6",
X"00000218",
X"000002e6",
X"00000118",
X"000000e6",
X"00000318",
X"00000366",
X"00000098",
X"00000166",
X"00000298",
X"00000266",
X"00000198",
X"00000066",
X"00000398",
X"000003a6",
X"00000058",
X"000001a6",
X"00000258",
X"000002a6",
X"00000158",
X"000000a6",
X"00000358",
X"00000326",
X"000000d8",
X"00000126",
X"000002d8",
X"00000226",
X"000001d8",
X"00000026",
X"000003d8",
X"000003c6",
X"00000038",
X"000001c6",
X"00000238",
X"000002c6",
X"00000138",
X"000000c6",
X"00000338",
X"00000346",
X"000000b8",
X"00000146",
X"000002b8",
X"00000246",
X"000001b8",
X"00000046",
X"000003b8",
X"00000386",
X"00000078",
X"00000186",
X"00000278",
X"00000286",
X"00000178",
X"00000086",
X"00000378",
X"00000306",
X"000000f8",
X"00000106",
X"000002f8",
X"00000206",
X"000001f8",
X"00000006",
X"000003f8",
X"000003fa",
X"00000004",
X"000001fa",
X"00000204",
X"000002fa",
X"00000104",
X"000000fa",
X"00000304",
X"0000037a",
X"00000084",
X"0000017a",
X"00000284",
X"0000027a",
X"00000184",
X"0000007a",
X"00000384",
X"000003ba",
X"00000044",
X"000001ba",
X"00000244",
X"000002ba",
X"00000144",
X"000000ba",
X"00000344",
X"0000033a",
X"000000c4",
X"0000013a",
X"000002c4",
X"0000023a",
X"000001c4",
X"0000003a",
X"000003c4",
X"000003da",
X"00000024",
X"000001da",
X"00000224",
X"000002da",
X"00000124",
X"000000da",
X"00000324",
X"0000035a",
X"000000a4",
X"0000015a",
X"000002a4",
X"0000025a",
X"000001a4",
X"0000005a",
X"000003a4",
X"0000039a",
X"00000064",
X"0000019a",
X"00000264",
X"0000029a",
X"00000164",
X"0000009a",
X"00000364",
X"0000031a",
X"000000e4",
X"0000011a",
X"000002e4",
X"0000021a",
X"000001e4",
X"0000001a",
X"000003e4",
X"000003ea",
X"00000014",
X"000001ea",
X"00000214",
X"000002ea",
X"00000114",
X"000000ea",
X"00000314",
X"0000036a",
X"00000094",
X"0000016a",
X"00000294",
X"0000026a",
X"00000194",
X"0000006a",
X"00000394",
X"000003aa",
X"00000054",
X"000001aa",
X"00000254",
X"000002aa",
X"00000154",
X"000000aa",
X"00000354",
X"0000032a",
X"000000d4",
X"0000012a",
X"000002d4",
X"0000022a",
X"000001d4",
X"0000002a",
X"000003d4",
X"000003ca",
X"00000034",
X"000001ca",
X"00000234",
X"000002ca",
X"00000134",
X"000000ca",
X"00000334",
X"0000034a",
X"000000b4",
X"0000014a",
X"000002b4",
X"0000024a",
X"000001b4",
X"0000004a",
X"000003b4",
X"0000038a",
X"00000074",
X"0000018a",
X"00000274",
X"0000028a",
X"00000174",
X"0000008a",
X"00000374",
X"0000030a",
X"000000f4",
X"0000010a",
X"000002f4",
X"0000020a",
X"000001f4",
X"0000000a",
X"000003f4",
X"000003f2",
X"0000000c",
X"000001f2",
X"0000020c",
X"000002f2",
X"0000010c",
X"000000f2",
X"0000030c",
X"00000372",
X"0000008c",
X"00000172",
X"0000028c",
X"00000272",
X"0000018c",
X"00000072",
X"0000038c",
X"000003b2",
X"0000004c",
X"000001b2",
X"0000024c",
X"000002b2",
X"0000014c",
X"000000b2",
X"0000034c",
X"00000332",
X"000000cc",
X"00000132",
X"000002cc",
X"00000232",
X"000001cc",
X"00000032",
X"000003cc",
X"000003d2",
X"0000002c",
X"000001d2",
X"0000022c",
X"000002d2",
X"0000012c",
X"000000d2",
X"0000032c",
X"00000352",
X"000000ac",
X"00000152",
X"000002ac",
X"00000252",
X"000001ac",
X"00000052",
X"000003ac",
X"00000392",
X"0000006c",
X"00000192",
X"0000026c",
X"00000292",
X"0000016c",
X"00000092",
X"0000036c",
X"00000312",
X"000000ec",
X"00000112",
X"000002ec",
X"00000212",
X"000001ec",
X"00000012",
X"000003ec",
X"000003e2",
X"0000001c",
X"000001e2",
X"0000021c",
X"000002e2",
X"0000011c",
X"000000e2",
X"0000031c",
X"00000362",
X"0000009c",
X"00000162",
X"0000029c",
X"00000262",
X"0000019c",
X"00000062",
X"0000039c",
X"000003a2",
X"0000005c",
X"000001a2",
X"0000025c",
X"000002a2",
X"0000015c",
X"000000a2",
X"0000035c",
X"00000322",
X"000000dc",
X"00000122",
X"000002dc",
X"00000222",
X"000001dc",
X"00000022",
X"000003dc",
X"000003c2",
X"0000003c",
X"000001c2",
X"0000023c",
X"000002c2",
X"0000013c",
X"000000c2",
X"0000033c",
X"00000342",
X"000000bc",
X"00000142",
X"000002bc",
X"00000242",
X"000001bc",
X"00000042",
X"000003bc",
X"00000382",
X"0000007c",
X"00000182",
X"0000027c",
X"00000282",
X"0000017c",
X"00000082",
X"0000037c",
X"00000302",
X"000000fc",
X"00000102",
X"000002fc",
X"00000202",
X"000001fc",
X"00000002",
X"000003fc"
);
--T:
constant T: rom_table:= rom_table'(
X"00004000",
X"00000000",
X"00003ffe",
X"ffffff9c",
X"00003ffd",
X"ffffff37",
X"00003ffc",
X"fffffed3",
X"00003ffb",
X"fffffe6e",
X"00003ff7",
X"fffffe0a",
X"00003ff3",
X"fffffda5",
X"00003fef",
X"fffffd41",
X"00003fec",
X"fffffcdc",
X"00003fe6",
X"fffffc78",
X"00003fe0",
X"fffffc14",
X"00003fda",
X"fffffbb0",
X"00003fd4",
X"fffffb4b",
X"00003fcb",
X"fffffae7",
X"00003fc2",
X"fffffa83",
X"00003fb9",
X"fffffa1f",
X"00003fb1",
X"fffff9ba",
X"00003fa6",
X"fffff956",
X"00003f9b",
X"fffff8f2",
X"00003f90",
X"fffff88e",
X"00003f85",
X"fffff82a",
X"00003f77",
X"fffff7c7",
X"00003f6a",
X"fffff763",
X"00003f5c",
X"fffff700",
X"00003f4f",
X"fffff69c",
X"00003f3f",
X"fffff639",
X"00003f2f",
X"fffff5d6",
X"00003f1f",
X"fffff573",
X"00003f0f",
X"fffff50f",
X"00003efc",
X"fffff4ad",
X"00003eea",
X"fffff44a",
X"00003ed7",
X"fffff3e7",
X"00003ec5",
X"fffff384",
X"00003eb0",
X"fffff322",
X"00003e9b",
X"fffff2bf",
X"00003e86",
X"fffff25d",
X"00003e72",
X"fffff1fa",
X"00003e5a",
X"fffff199",
X"00003e43",
X"fffff137",
X"00003e2c",
X"fffff0d5",
X"00003e15",
X"fffff073",
X"00003dfb",
X"fffff012",
X"00003de2",
X"ffffefb1",
X"00003dc8",
X"ffffef50",
X"00003daf",
X"ffffeeee",
X"00003d93",
X"ffffee8e",
X"00003d77",
X"ffffee2d",
X"00003d5b",
X"ffffedcd",
X"00003d3f",
X"ffffed6c",
X"00003d20",
X"ffffed0d",
X"00003d02",
X"ffffecad",
X"00003ce3",
X"ffffec4d",
X"00003cc5",
X"ffffebed",
X"00003ca4",
X"ffffeb8e",
X"00003c83",
X"ffffeb2f",
X"00003c62",
X"ffffead0",
X"00003c42",
X"ffffea70",
X"00003c1f",
X"ffffea12",
X"00003bfc",
X"ffffe9b4",
X"00003bd9",
X"ffffe956",
X"00003bb6",
X"ffffe8f7",
X"00003b90",
X"ffffe89a",
X"00003b6b",
X"ffffe83d",
X"00003b46",
X"ffffe7e0",
X"00003b21",
X"ffffe782",
X"00003af9",
X"ffffe726",
X"00003ad1",
X"ffffe6ca",
X"00003aa9",
X"ffffe66e",
X"00003a82",
X"ffffe611",
X"00003a58",
X"ffffe5b6",
X"00003a2e",
X"ffffe55a",
X"00003a04",
X"ffffe4ff",
X"000039db",
X"ffffe4a3",
X"000039af",
X"ffffe449",
X"00003983",
X"ffffe3ef",
X"00003957",
X"ffffe395",
X"0000392b",
X"ffffe33a",
X"000038fc",
X"ffffe2e1",
X"000038ce",
X"ffffe288",
X"0000389f",
X"ffffe22f",
X"00003871",
X"ffffe1d5",
X"00003840",
X"ffffe17d",
X"00003810",
X"ffffe125",
X"000037e0",
X"ffffe0cd",
X"000037b0",
X"ffffe074",
X"0000377d",
X"ffffe01e",
X"0000374a",
X"ffffdfc7",
X"00003717",
X"ffffdf70",
X"000036e5",
X"ffffdf19",
X"000036b0",
X"ffffdec4",
X"0000367b",
X"ffffde6e",
X"00003646",
X"ffffde19",
X"00003612",
X"ffffddc3",
X"000035db",
X"ffffdd6f",
X"000035a4",
X"ffffdd1b",
X"0000356d",
X"ffffdcc7",
X"00003537",
X"ffffdc72",
X"000034fe",
X"ffffdc1f",
X"000034c5",
X"ffffdbcc",
X"0000348c",
X"ffffdb79",
X"00003453",
X"ffffdb26",
X"00003418",
X"ffffdad5",
X"000033dd",
X"ffffda83",
X"000033a2",
X"ffffda32",
X"00003368",
X"ffffd9e0",
X"0000332b",
X"ffffd990",
X"000032ee",
X"ffffd940",
X"000032b1",
X"ffffd8f0",
X"00003274",
X"ffffd8a0",
X"00003235",
X"ffffd852",
X"000031f6",
X"ffffd803",
X"000031b7",
X"ffffd7b5",
X"00003179",
X"ffffd766",
X"00003138",
X"ffffd719",
X"000030f7",
X"ffffd6cc",
X"000030b6",
X"ffffd67f",
X"00003076",
X"ffffd632",
X"00003033",
X"ffffd5e7",
X"00002ff1",
X"ffffd59c",
X"00002fae",
X"ffffd551",
X"00002f6c",
X"ffffd505",
X"00002f27",
X"ffffd4bc",
X"00002ee3",
X"ffffd472",
X"00002e9e",
X"ffffd429",
X"00002e5a",
X"ffffd3df",
X"00002e13",
X"ffffd397",
X"00002dcd",
X"ffffd34f",
X"00002d87",
X"ffffd307",
X"00002d41",
X"ffffd2bf",
X"00002cf9",
X"ffffd279",
X"00002cb1",
X"ffffd233",
X"00002c69",
X"ffffd1ed",
X"00002c21",
X"ffffd1a6",
X"00002bd7",
X"ffffd162",
X"00002b8e",
X"ffffd11d",
X"00002b44",
X"ffffd0d9",
X"00002afb",
X"ffffd094",
X"00002aaf",
X"ffffd052",
X"00002a64",
X"ffffd00f",
X"00002a19",
X"ffffcfcd",
X"000029ce",
X"ffffcf8a",
X"00002981",
X"ffffcf4a",
X"00002934",
X"ffffcf09",
X"000028e7",
X"ffffcec8",
X"0000289a",
X"ffffce87",
X"0000284b",
X"ffffce49",
X"000027fd",
X"ffffce0a",
X"000027ae",
X"ffffcdcb",
X"00002760",
X"ffffcd8c",
X"00002710",
X"ffffcd4f",
X"000026c0",
X"ffffcd12",
X"00002670",
X"ffffccd5",
X"00002620",
X"ffffcc98",
X"000025ce",
X"ffffcc5e",
X"0000257d",
X"ffffcc23",
X"0000252b",
X"ffffcbe8",
X"000024da",
X"ffffcbad",
X"00002487",
X"ffffcb74",
X"00002434",
X"ffffcb3b",
X"000023e1",
X"ffffcb02",
X"0000238e",
X"ffffcac9",
X"00002339",
X"ffffca93",
X"000022e5",
X"ffffca5c",
X"00002291",
X"ffffca25",
X"0000223d",
X"ffffc9ee",
X"000021e7",
X"ffffc9ba",
X"00002192",
X"ffffc985",
X"0000213c",
X"ffffc950",
X"000020e7",
X"ffffc91b",
X"00002090",
X"ffffc8e9",
X"00002039",
X"ffffc8b6",
X"00001fe2",
X"ffffc883",
X"00001f8c",
X"ffffc850",
X"00001f33",
X"ffffc820",
X"00001edb",
X"ffffc7f0",
X"00001e83",
X"ffffc7c0",
X"00001e2b",
X"ffffc78f",
X"00001dd1",
X"ffffc761",
X"00001d78",
X"ffffc732",
X"00001d1f",
X"ffffc704",
X"00001cc6",
X"ffffc6d5",
X"00001c6b",
X"ffffc6a9",
X"00001c11",
X"ffffc67d",
X"00001bb7",
X"ffffc651",
X"00001b5d",
X"ffffc625",
X"00001b01",
X"ffffc5fc",
X"00001aa6",
X"ffffc5d2",
X"00001a4a",
X"ffffc5a8",
X"000019ef",
X"ffffc57e",
X"00001992",
X"ffffc557",
X"00001936",
X"ffffc52f",
X"000018da",
X"ffffc507",
X"0000187e",
X"ffffc4df",
X"00001820",
X"ffffc4ba",
X"000017c3",
X"ffffc495",
X"00001766",
X"ffffc470",
X"00001709",
X"ffffc44a",
X"000016aa",
X"ffffc427",
X"0000164c",
X"ffffc404",
X"000015ee",
X"ffffc3e1",
X"00001590",
X"ffffc3be",
X"00001530",
X"ffffc39e",
X"000014d1",
X"ffffc37d",
X"00001472",
X"ffffc35c",
X"00001413",
X"ffffc33b",
X"000013b3",
X"ffffc31d",
X"00001353",
X"ffffc2fe",
X"000012f3",
X"ffffc2e0",
X"00001294",
X"ffffc2c1",
X"00001233",
X"ffffc2a5",
X"000011d3",
X"ffffc289",
X"00001172",
X"ffffc26d",
X"00001112",
X"ffffc251",
X"000010b0",
X"ffffc238",
X"0000104f",
X"ffffc21e",
X"00000fee",
X"ffffc205",
X"00000f8d",
X"ffffc1eb",
X"00000f2b",
X"ffffc1d4",
X"00000ec9",
X"ffffc1bd",
X"00000e67",
X"ffffc1a6",
X"00000e06",
X"ffffc18e",
X"00000da3",
X"ffffc17a",
X"00000d41",
X"ffffc165",
X"00000cde",
X"ffffc150",
X"00000c7c",
X"ffffc13b",
X"00000c19",
X"ffffc129",
X"00000bb6",
X"ffffc116",
X"00000b53",
X"ffffc104",
X"00000af1",
X"ffffc0f1",
X"00000a8d",
X"ffffc0e1",
X"00000a2a",
X"ffffc0d1",
X"000009c7",
X"ffffc0c1",
X"00000964",
X"ffffc0b1",
X"00000900",
X"ffffc0a4",
X"0000089d",
X"ffffc096",
X"00000839",
X"ffffc089",
X"000007d6",
X"ffffc07b",
X"00000772",
X"ffffc070",
X"0000070e",
X"ffffc065",
X"000006aa",
X"ffffc05a",
X"00000646",
X"ffffc04f",
X"000005e1",
X"ffffc047",
X"0000057d",
X"ffffc03e",
X"00000519",
X"ffffc035",
X"000004b5",
X"ffffc02c",
X"00000450",
X"ffffc026",
X"000003ec",
X"ffffc020",
X"00000388",
X"ffffc01a",
X"00000324",
X"ffffc014",
X"000002bf",
X"ffffc011",
X"0000025b",
X"ffffc00d",
X"000001f6",
X"ffffc009",
X"00000192",
X"ffffc005",
X"0000012d",
X"ffffc004",
X"000000c9",
X"ffffc003",
X"00000064",
X"ffffc002",
X"00000000",
X"ffffc000",
X"ffffff9b",
X"ffffc002",
X"ffffff37",
X"ffffc003",
X"fffffed3",
X"ffffc004",
X"fffffe6f",
X"ffffc005",
X"fffffe0a",
X"ffffc009",
X"fffffda6",
X"ffffc00d",
X"fffffd41",
X"ffffc011",
X"fffffcdd",
X"ffffc014",
X"fffffc78",
X"ffffc01a",
X"fffffc14",
X"ffffc020",
X"fffffbb0",
X"ffffc026",
X"fffffb4c",
X"ffffc02c",
X"fffffae7",
X"ffffc035",
X"fffffa83",
X"ffffc03e",
X"fffffa1f",
X"ffffc047",
X"fffff9bb",
X"ffffc04f",
X"fffff957",
X"ffffc05a",
X"fffff8f3",
X"ffffc065",
X"fffff88f",
X"ffffc070",
X"fffff82b",
X"ffffc07b",
X"fffff7c7",
X"ffffc089",
X"fffff764",
X"ffffc096",
X"fffff700",
X"ffffc0a4",
X"fffff69d",
X"ffffc0b1",
X"fffff639",
X"ffffc0c1",
X"fffff5d6",
X"ffffc0d1",
X"fffff573",
X"ffffc0e1",
X"fffff510",
X"ffffc0f1",
X"fffff4ad",
X"ffffc104",
X"fffff44a",
X"ffffc116",
X"fffff3e7",
X"ffffc129",
X"fffff385",
X"ffffc13b",
X"fffff322",
X"ffffc150",
X"fffff2c0",
X"ffffc165",
X"fffff25d",
X"ffffc17a",
X"fffff1fb",
X"ffffc18e",
X"fffff199",
X"ffffc1a6",
X"fffff137",
X"ffffc1bd",
X"fffff0d5",
X"ffffc1d4",
X"fffff074",
X"ffffc1eb",
X"fffff012",
X"ffffc205",
X"ffffefb1",
X"ffffc21e",
X"ffffef50",
X"ffffc238",
X"ffffeeef",
X"ffffc251",
X"ffffee8e",
X"ffffc26d",
X"ffffee2e",
X"ffffc289",
X"ffffedcd",
X"ffffc2a5",
X"ffffed6d",
X"ffffc2c1",
X"ffffed0d",
X"ffffc2e0",
X"ffffecad",
X"ffffc2fe",
X"ffffec4d",
X"ffffc31d",
X"ffffebee",
X"ffffc33b",
X"ffffeb8e",
X"ffffc35c",
X"ffffeb2f",
X"ffffc37d",
X"ffffead0",
X"ffffc39e",
X"ffffea71",
X"ffffc3be",
X"ffffea12",
X"ffffc3e1",
X"ffffe9b4",
X"ffffc404",
X"ffffe956",
X"ffffc427",
X"ffffe8f8",
X"ffffc44a",
X"ffffe89a",
X"ffffc470",
X"ffffe83d",
X"ffffc495",
X"ffffe7e0",
X"ffffc4ba",
X"ffffe783",
X"ffffc4df",
X"ffffe726",
X"ffffc507",
X"ffffe6ca",
X"ffffc52f",
X"ffffe66e",
X"ffffc557",
X"ffffe612",
X"ffffc57e",
X"ffffe5b6",
X"ffffc5a8",
X"ffffe55b",
X"ffffc5d2",
X"ffffe4ff",
X"ffffc5fc",
X"ffffe4a4",
X"ffffc625",
X"ffffe449",
X"ffffc651",
X"ffffe3ef",
X"ffffc67d",
X"ffffe395",
X"ffffc6a9",
X"ffffe33b",
X"ffffc6d5",
X"ffffe2e1",
X"ffffc704",
X"ffffe288",
X"ffffc732",
X"ffffe22f",
X"ffffc761",
X"ffffe1d6",
X"ffffc78f",
X"ffffe17d",
X"ffffc7c0",
X"ffffe125",
X"ffffc7f0",
X"ffffe0cd",
X"ffffc820",
X"ffffe075",
X"ffffc850",
X"ffffe01e",
X"ffffc883",
X"ffffdfc7",
X"ffffc8b6",
X"ffffdf70",
X"ffffc8e9",
X"ffffdf1a",
X"ffffc91b",
X"ffffdec4",
X"ffffc950",
X"ffffde6f",
X"ffffc985",
X"ffffde19",
X"ffffc9ba",
X"ffffddc4",
X"ffffc9ee",
X"ffffdd6f",
X"ffffca25",
X"ffffdd1b",
X"ffffca5c",
X"ffffdcc7",
X"ffffca93",
X"ffffdc73",
X"ffffcac9",
X"ffffdc20",
X"ffffcb02",
X"ffffdbcd",
X"ffffcb3b",
X"ffffdb7a",
X"ffffcb74",
X"ffffdb27",
X"ffffcbad",
X"ffffdad5",
X"ffffcbe8",
X"ffffda84",
X"ffffcc23",
X"ffffda32",
X"ffffcc5e",
X"ffffd9e1",
X"ffffcc98",
X"ffffd991",
X"ffffccd5",
X"ffffd941",
X"ffffcd12",
X"ffffd8f1",
X"ffffcd4f",
X"ffffd8a1",
X"ffffcd8c",
X"ffffd852",
X"ffffcdcb",
X"ffffd804",
X"ffffce0a",
X"ffffd7b5",
X"ffffce49",
X"ffffd767",
X"ffffce87",
X"ffffd71a",
X"ffffcec8",
X"ffffd6cd",
X"ffffcf09",
X"ffffd680",
X"ffffcf4a",
X"ffffd633",
X"ffffcf8a",
X"ffffd5e7",
X"ffffcfcd",
X"ffffd59c",
X"ffffd00f",
X"ffffd551",
X"ffffd052",
X"ffffd506",
X"ffffd094",
X"ffffd4bc",
X"ffffd0d9",
X"ffffd473",
X"ffffd11d",
X"ffffd429",
X"ffffd162",
X"ffffd3e0",
X"ffffd1a6",
X"ffffd398",
X"ffffd1ed",
X"ffffd350",
X"ffffd233",
X"ffffd308",
X"ffffd279",
X"ffffd2c0",
X"ffffd2bf",
X"ffffd279",
X"ffffd307",
X"ffffd233",
X"ffffd34f",
X"ffffd1ed",
X"ffffd397",
X"ffffd1a7",
X"ffffd3df",
X"ffffd162",
X"ffffd429",
X"ffffd11e",
X"ffffd472",
X"ffffd0d9",
X"ffffd4bc",
X"ffffd095",
X"ffffd505",
X"ffffd052",
X"ffffd551",
X"ffffd010",
X"ffffd59c",
X"ffffcfcd",
X"ffffd5e7",
X"ffffcf8b",
X"ffffd632",
X"ffffcf4a",
X"ffffd67f",
X"ffffcf09",
X"ffffd6cc",
X"ffffcec8",
X"ffffd719",
X"ffffce88",
X"ffffd766",
X"ffffce49",
X"ffffd7b5",
X"ffffce0a",
X"ffffd803",
X"ffffcdcb",
X"ffffd852",
X"ffffcd8d",
X"ffffd8a0",
X"ffffcd50",
X"ffffd8f0",
X"ffffcd13",
X"ffffd940",
X"ffffccd6",
X"ffffd990",
X"ffffcc99",
X"ffffd9e0",
X"ffffcc5e",
X"ffffda32",
X"ffffcc23",
X"ffffda83",
X"ffffcbe8",
X"ffffdad5",
X"ffffcbae",
X"ffffdb26",
X"ffffcb75",
X"ffffdb79",
X"ffffcb3c",
X"ffffdbcc",
X"ffffcb03",
X"ffffdc1f",
X"ffffcaca",
X"ffffdc72",
X"ffffca93",
X"ffffdcc7",
X"ffffca5c",
X"ffffdd1b",
X"ffffca25",
X"ffffdd6f",
X"ffffc9ef",
X"ffffddc3",
X"ffffc9ba",
X"ffffde19",
X"ffffc985",
X"ffffde6e",
X"ffffc950",
X"ffffdec4",
X"ffffc91c",
X"ffffdf19",
X"ffffc8e9",
X"ffffdf70",
X"ffffc8b6",
X"ffffdfc7",
X"ffffc883",
X"ffffe01e",
X"ffffc851",
X"ffffe074",
X"ffffc820",
X"ffffe0cd",
X"ffffc7f0",
X"ffffe125",
X"ffffc7c0",
X"ffffe17d",
X"ffffc790",
X"ffffe1d5",
X"ffffc761",
X"ffffe22f",
X"ffffc733",
X"ffffe288",
X"ffffc704",
X"ffffe2e1",
X"ffffc6d6",
X"ffffe33a",
X"ffffc6aa",
X"ffffe395",
X"ffffc67e",
X"ffffe3ef",
X"ffffc652",
X"ffffe449",
X"ffffc626",
X"ffffe4a3",
X"ffffc5fc",
X"ffffe4ff",
X"ffffc5d2",
X"ffffe55a",
X"ffffc5a8",
X"ffffe5b6",
X"ffffc57f",
X"ffffe611",
X"ffffc557",
X"ffffe66e",
X"ffffc52f",
X"ffffe6ca",
X"ffffc507",
X"ffffe726",
X"ffffc4e0",
X"ffffe782",
X"ffffc4ba",
X"ffffe7e0",
X"ffffc495",
X"ffffe83d",
X"ffffc470",
X"ffffe89a",
X"ffffc44b",
X"ffffe8f7",
X"ffffc428",
X"ffffe956",
X"ffffc405",
X"ffffe9b4",
X"ffffc3e2",
X"ffffea12",
X"ffffc3bf",
X"ffffea70",
X"ffffc39e",
X"ffffead0",
X"ffffc37d",
X"ffffeb2f",
X"ffffc35c",
X"ffffeb8e",
X"ffffc33c",
X"ffffebed",
X"ffffc31d",
X"ffffec4d",
X"ffffc2ff",
X"ffffecad",
X"ffffc2e0",
X"ffffed0d",
X"ffffc2c2",
X"ffffed6c",
X"ffffc2a6",
X"ffffedcd",
X"ffffc28a",
X"ffffee2d",
X"ffffc26e",
X"ffffee8e",
X"ffffc252",
X"ffffeeee",
X"ffffc238",
X"ffffef50",
X"ffffc21f",
X"ffffefb1",
X"ffffc205",
X"fffff012",
X"ffffc1ec",
X"fffff073",
X"ffffc1d4",
X"fffff0d5",
X"ffffc1bd",
X"fffff137",
X"ffffc1a6",
X"fffff199",
X"ffffc18f",
X"fffff1fa",
X"ffffc17a",
X"fffff25d",
X"ffffc165",
X"fffff2bf",
X"ffffc150",
X"fffff322",
X"ffffc13c",
X"fffff384",
X"ffffc129",
X"fffff3e7",
X"ffffc117",
X"fffff44a",
X"ffffc104",
X"fffff4ad",
X"ffffc0f2",
X"fffff50f",
X"ffffc0e2",
X"fffff573",
X"ffffc0d2",
X"fffff5d6",
X"ffffc0c2",
X"fffff639",
X"ffffc0b2",
X"fffff69c",
X"ffffc0a4",
X"fffff700",
X"ffffc097",
X"fffff763",
X"ffffc089",
X"fffff7c7",
X"ffffc07c",
X"fffff82a",
X"ffffc071",
X"fffff88e",
X"ffffc066",
X"fffff8f2",
X"ffffc05b",
X"fffff956",
X"ffffc050",
X"fffff9ba",
X"ffffc047",
X"fffffa1f",
X"ffffc03e",
X"fffffa83",
X"ffffc035",
X"fffffae7",
X"ffffc02d",
X"fffffb4b",
X"ffffc027",
X"fffffbb0",
X"ffffc021",
X"fffffc14",
X"ffffc01b",
X"fffffc78",
X"ffffc015",
X"fffffcdc",
X"ffffc011",
X"fffffd41",
X"ffffc00d",
X"fffffda5",
X"ffffc009",
X"fffffe0a",
X"ffffc006",
X"fffffe6e",
X"ffffc004",
X"fffffed3",
X"ffffc003",
X"ffffff37",
X"ffffc002",
X"ffffff9c",
X"00003fff",
X"0000000c",
X"00003fff",
X"00000025",
X"00003fff",
X"0000003e",
X"00003ffe",
X"00000057",
X"00003ffe",
X"00000071",
X"00003ffe",
X"0000008a",
X"00003ffd",
X"000000a3",
X"00003ffd",
X"000000bc",
X"00003ffd",
X"000000d5",
X"00003ffd",
X"000000ee",
X"00003ffc",
X"00000107",
X"00003ffc",
X"00000120",
X"00003ffc",
X"0000013a",
X"00003ffb",
X"00000153",
X"00003ffb",
X"0000016c",
X"00003ffb",
X"00000185",
X"00003ffa",
X"0000019e",
X"00003ff9",
X"000001b7",
X"00003ff8",
X"000001d0",
X"00003ff7",
X"000001e9",
X"00003ff6",
X"00000203",
X"00003ff5",
X"0000021c",
X"00003ff4",
X"00000235",
X"00003ff3",
X"0000024e",
X"00003ff3",
X"00000267",
X"00003ff2",
X"00000280",
X"00003ff1",
X"00000299",
X"00003ff0",
X"000002b2",
X"00003fef",
X"000002cc",
X"00003fee",
X"000002e5",
X"00003fed",
X"000002fe",
X"00003fec",
X"00000317",
X"00003feb",
X"00000330",
X"00003fe9",
X"00000349",
X"00003fe8",
X"00000362",
X"00003fe6",
X"0000037b",
X"00003fe5",
X"00000394",
X"00003fe3",
X"000003ad",
X"00003fe2",
X"000003c6",
X"00003fe0",
X"000003df",
X"00003fdf",
X"000003f9",
X"00003fdd",
X"00000412",
X"00003fdc",
X"0000042b",
X"00003fda",
X"00000444",
X"00003fd9",
X"0000045d",
X"00003fd7",
X"00000476",
X"00003fd6",
X"0000048f",
X"00003fd4",
X"000004a8",
X"00003fd2",
X"000004c1",
X"00003fd0",
X"000004da",
X"00003fce",
X"000004f3",
X"00003fcc",
X"0000050c",
X"00003fca",
X"00000525",
X"00003fc7",
X"0000053e",
X"00003fc5",
X"00000557",
X"00003fc3",
X"00000570",
X"00003fc1",
X"0000058a",
X"00003fbf",
X"000005a3",
X"00003fbd",
X"000005bc",
X"00003fba",
X"000005d5",
X"00003fb8",
X"000005ee",
X"00003fb6",
X"00000607",
X"00003fb4",
X"00000620",
X"00003fb2",
X"00000639",
X"00003faf",
X"00000652",
X"00003fac",
X"0000066b",
X"00003faa",
X"00000684",
X"00003fa7",
X"0000069d",
X"00003fa4",
X"000006b6",
X"00003fa1",
X"000006cf",
X"00003f9f",
X"000006e8",
X"00003f9c",
X"00000701",
X"00003f99",
X"0000071a",
X"00003f96",
X"00000733",
X"00003f94",
X"0000074c",
X"00003f91",
X"00000765",
X"00003f8e",
X"0000077e",
X"00003f8b",
X"00000797",
X"00003f89",
X"000007b0",
X"00003f86",
X"000007c9",
X"00003f83",
X"000007e2",
X"00003f7f",
X"000007fb",
X"00003f7c",
X"00000814",
X"00003f79",
X"0000082d",
X"00003f75",
X"00000845",
X"00003f72",
X"0000085e",
X"00003f6f",
X"00000877",
X"00003f6b",
X"00000890",
X"00003f68",
X"000008a9",
X"00003f64",
X"000008c2",
X"00003f61",
X"000008db",
X"00003f5e",
X"000008f4",
X"00003f5a",
X"0000090c",
X"00003f57",
X"00000925",
X"00003f54",
X"0000093e",
X"00003f50",
X"00000957",
X"00003f4d",
X"00000970",
X"00003f49",
X"00000989",
X"00003f45",
X"000009a2",
X"00003f41",
X"000009ba",
X"00003f3d",
X"000009d3",
X"00003f39",
X"000009ec",
X"00003f35",
X"00000a05",
X"00003f31",
X"00000a1e",
X"00003f2d",
X"00000a36",
X"00003f29",
X"00000a4f",
X"00003f25",
X"00000a68",
X"00003f21",
X"00000a81",
X"00003f1d",
X"00000a9a",
X"00003f19",
X"00000ab2",
X"00003f15",
X"00000acb",
X"00003f11",
X"00000ae4",
X"00003f0c",
X"00000afd",
X"00003f08",
X"00000b16",
X"00003f03",
X"00000b2e",
X"00003efe",
X"00000b47",
X"00003efa",
X"00000b60",
X"00003ef5",
X"00000b78",
X"00003ef0",
X"00000b91",
X"00003eec",
X"00000baa",
X"00003ee7",
X"00000bc2",
X"00003ee3",
X"00000bdb",
X"00003ede",
X"00000bf4",
X"00003ed9",
X"00000c0c",
X"00003ed5",
X"00000c25",
X"00003ed0",
X"00000c3e",
X"00003ecb",
X"00000c56",
X"00003ec7",
X"00000c6f",
X"00003ec2",
X"00000c88",
X"00003ebd",
X"00000ca0",
X"00003eb8",
X"00000cb9",
X"00003eb2",
X"00000cd2",
X"00003ead",
X"00000cea",
X"00003ea8",
X"00000d03",
X"00003ea3",
X"00000d1c",
X"00003e9e",
X"00000d34",
X"00003e98",
X"00000d4d",
X"00003e93",
X"00000d65",
X"00003e8e",
X"00000d7e",
X"00003e89",
X"00000d97",
X"00003e84",
X"00000daf",
X"00003e7e",
X"00000dc8",
X"00003e79",
X"00000de1",
X"00003e74",
X"00000df9",
X"00003e6f",
X"00000e12",
X"00003e69",
X"00000e2a",
X"00003e63",
X"00000e43",
X"00003e5d",
X"00000e5b",
X"00003e57",
X"00000e73",
X"00003e52",
X"00000e8c",
X"00003e4c",
X"00000ea4",
X"00003e46",
X"00000ebd",
X"00003e40",
X"00000ed5",
X"00003e3a",
X"00000eee",
X"00003e34",
X"00000f06",
X"00003e2f",
X"00000f1f",
X"00003e29",
X"00000f37",
X"00003e23",
X"00000f4f",
X"00003e1d",
X"00000f68",
X"00003e17",
X"00000f80",
X"00003e11",
X"00000f99",
X"00003e0b",
X"00000fb1",
X"00003e05",
X"00000fc9",
X"00003dfe",
X"00000fe2",
X"00003df8",
X"00000ffa",
X"00003df1",
X"00001012",
X"00003deb",
X"0000102b",
X"00003de5",
X"00001043",
X"00003dde",
X"0000105b",
X"00003dd8",
X"00001073",
X"00003dd2",
X"0000108c",
X"00003dcb",
X"000010a4",
X"00003dc5",
X"000010bc",
X"00003dbe",
X"000010d5",
X"00003db8",
X"000010ed",
X"00003db2",
X"00001105",
X"00003dab",
X"0000111e",
X"00003da4",
X"00001136",
X"00003d9d",
X"0000114e",
X"00003d96",
X"00001166",
X"00003d8f",
X"0000117e",
X"00003d88",
X"00001196",
X"00003d81",
X"000011ae",
X"00003d7a",
X"000011c6",
X"00003d73",
X"000011df",
X"00003d6c",
X"000011f7",
X"00003d65",
X"0000120f",
X"00003d5e",
X"00001227",
X"00003d57",
X"0000123f",
X"00003d50",
X"00001257",
X"00003d49",
X"0000126f",
X"00003d42",
X"00001287",
X"00003d3b",
X"0000129f",
X"00003d33",
X"000012b7",
X"00003d2b",
X"000012cf",
X"00003d24",
X"000012e7",
X"00003d1c",
X"000012ff",
X"00003d15",
X"00001317",
X"00003d0d",
X"0000132f",
X"00003d05",
X"00001347",
X"00003cfe",
X"0000135f",
X"00003cf6",
X"00001377",
X"00003cee",
X"0000138f",
X"00003ce7",
X"000013a7",
X"00003cdf",
X"000013bf",
X"00003cd8",
X"000013d7",
X"00003cd0",
X"000013ef",
X"00003cc8",
X"00001407",
X"00003cc0",
X"0000141e",
X"00003cb8",
X"00001436",
X"00003cb0",
X"0000144e",
X"00003ca8",
X"00001466",
X"00003ca0",
X"0000147e",
X"00003c97",
X"00001495",
X"00003c8f",
X"000014ad",
X"00003c87",
X"000014c5",
X"00003c7f",
X"000014dd",
X"00003c77",
X"000014f5",
X"00003c6f",
X"0000150d",
X"00003c66",
X"00001524",
X"00003c5e",
X"0000153c",
X"00003c56",
X"00001554",
X"00003c4e",
X"0000156c",
X"00003c46",
X"00001584",
X"00003c3d",
X"0000159b",
X"00003c34",
X"000015b3",
X"00003c2c",
X"000015ca",
X"00003c23",
X"000015e2",
X"00003c1a",
X"000015fa",
X"00003c11",
X"00001611",
X"00003c09",
X"00001629",
X"00003c00",
X"00001640",
X"00003bf7",
X"00001658",
X"00003bee",
X"0000166f",
X"00003be6",
X"00001687",
X"00003bdd",
X"0000169e",
X"00003bd4",
X"000016b6",
X"00003bcb",
X"000016ce",
X"00003bc3",
X"000016e5",
X"00003bba",
X"000016fd",
X"00003bb1",
X"00001714",
X"00003ba8",
X"0000172b",
X"00003b9e",
X"00001743",
X"00003b95",
X"0000175a",
X"00003b8c",
X"00001771",
X"00003b82",
X"00001789",
X"00003b79",
X"000017a0",
X"00003b70",
X"000017b7",
X"00003b66",
X"000017cf",
X"00003b5d",
X"000017e6",
X"00003b54",
X"000017fd",
X"00003b4a",
X"00001815",
X"00003b41",
X"0000182c",
X"00003b38",
X"00001843",
X"00003b2e",
X"0000185b",
X"00003b25",
X"00001872",
X"00003b1c",
X"00001889",
X"00003b12",
X"000018a0",
X"00003b08",
X"000018b7",
X"00003afe",
X"000018ce",
X"00003af4",
X"000018e5",
X"00003aea",
X"000018fc",
X"00003ae0",
X"00001913",
X"00003ad6",
X"0000192a",
X"00003acc",
X"00001942",
X"00003ac2",
X"00001959",
X"00003ab8",
X"00001970",
X"00003aae",
X"00001987",
X"00003aa4",
X"0000199e",
X"00003a9a",
X"000019b5",
X"00003a90",
X"000019cc",
X"00003a86",
X"000019e3",
X"00003a7c",
X"000019fa",
X"00003a72",
X"00001a11",
X"00003a67",
X"00001a28",
X"00003a5d",
X"00001a3f",
X"00003a53",
X"00001a55",
X"00003a48",
X"00001a6c",
X"00003a3e",
X"00001a83",
X"00003a33",
X"00001a9a",
X"00003a29",
X"00001ab1",
X"00003a1e",
X"00001ac8",
X"00003a14",
X"00001adf",
X"00003a09",
X"00001af6",
X"000039ff",
X"00001b0c",
X"000039f5",
X"00001b23",
X"000039ea",
X"00001b3a",
X"000039e0",
X"00001b51",
X"000039d5",
X"00001b68",
X"000039ca",
X"00001b7e",
X"000039bf",
X"00001b95",
X"000039b4",
X"00001bab",
X"000039a9",
X"00001bc2",
X"0000399e",
X"00001bd9",
X"00003993",
X"00001bef",
X"00003988",
X"00001c06",
X"0000397d",
X"00001c1c",
X"00003972",
X"00001c33",
X"00003967",
X"00001c49",
X"0000395c",
X"00001c60",
X"00003951",
X"00001c77",
X"00003946",
X"00001c8d",
X"0000393b",
X"00001ca4",
X"00003930",
X"00001cba",
X"00003925",
X"00001cd1",
X"00003919",
X"00001ce7",
X"0000390d",
X"00001cfd",
X"00003902",
X"00001d14",
X"000038f6",
X"00001d2a",
X"000038eb",
X"00001d40",
X"000038df",
X"00001d57",
X"000038d3",
X"00001d6d",
X"000038c8",
X"00001d83",
X"000038bc",
X"00001d99",
X"000038b0",
X"00001db0",
X"000038a5",
X"00001dc6",
X"00003899",
X"00001ddc",
X"0000388e",
X"00001df3",
X"00003882",
X"00001e09",
X"00003876",
X"00001e1f",
X"0000386a",
X"00001e36",
X"0000385e",
X"00001e4c",
X"00003852",
X"00001e62",
X"00003846",
X"00001e78",
X"0000383a",
X"00001e8e",
X"0000382e",
X"00001ea4",
X"00003822",
X"00001eba",
X"00003816",
X"00001ed0",
X"0000380a",
X"00001ee6",
X"000037fe",
X"00001efc",
X"000037f2",
X"00001f12",
X"000037e6",
X"00001f28",
X"000037da",
X"00001f3e",
X"000037ce",
X"00001f54",
X"000037c2",
X"00001f6a",
X"000037b6",
X"00001f80",
X"000037a9",
X"00001f96",
X"0000379c",
X"00001fac",
X"00003790",
X"00001fc2",
X"00003783",
X"00001fd7",
X"00003776",
X"00001fed",
X"0000376a",
X"00002003",
X"0000375d",
X"00002018",
X"00003750",
X"0000202e",
X"00003744",
X"00002044",
X"00003737",
X"0000205a",
X"0000372a",
X"0000206f",
X"0000371e",
X"00002085",
X"00003711",
X"0000209b",
X"00003704",
X"000020b0",
X"000036f8",
X"000020c6",
X"000036eb",
X"000020dc",
X"000036de",
X"000020f1",
X"000036d1",
X"00002107",
X"000036c4",
X"0000211c",
X"000036b6",
X"00002131",
X"000036a9",
X"00002147",
X"0000369c",
X"0000215c",
X"0000368f",
X"00002171",
X"00003682",
X"00002187",
X"00003674",
X"0000219c",
X"00003667",
X"000021b2",
X"0000365a",
X"000021c7",
X"0000364d",
X"000021dc",
X"00003640",
X"000021f2",
X"00003632",
X"00002207",
X"00003625",
X"0000221c",
X"00003618",
X"00002232",
X"0000360b",
X"00002247",
X"000035fd",
X"0000225c",
X"000035ef",
X"00002271",
X"000035e2",
X"00002286",
X"000035d4",
X"0000229b",
X"000035c6",
X"000022b0",
X"000035b9",
X"000022c5",
X"000035ab",
X"000022da",
X"0000359d",
X"000022f0",
X"0000358f",
X"00002305",
X"00003582",
X"0000231a",
X"00003574",
X"0000232f",
X"00003566",
X"00002344",
X"00003559",
X"00002359",
X"0000354b",
X"0000236e",
X"0000353d",
X"00002383",
X"0000352f",
X"00002398",
X"00003521",
X"000023ad",
X"00003513",
X"000023c1",
X"00003505",
X"000023d6",
X"000034f6",
X"000023eb",
X"000034e8",
X"00002400",
X"000034da",
X"00002414",
X"000034cc",
X"00002429",
X"000034bd",
X"0000243e",
X"000034af",
X"00002453",
X"000034a1",
X"00002467",
X"00003493",
X"0000247c",
X"00003484",
X"00002491",
X"00003476",
X"000024a6",
X"00003468",
X"000024ba",
X"0000345a",
X"000024cf",
X"0000344b",
X"000024e4",
X"0000343c",
X"000024f8",
X"0000342e",
X"0000250c",
X"0000341f",
X"00002521",
X"00003410",
X"00002535",
X"00003402",
X"0000254a",
X"000033f3",
X"0000255e",
X"000033e4",
X"00002572",
X"000033d6",
X"00002587",
X"000033c7",
X"0000259b",
X"000033b8",
X"000025af",
X"000033aa",
X"000025c4",
X"0000339b",
X"000025d8",
X"0000338c",
X"000025ed",
X"0000337e",
X"00002601",
X"0000336f",
X"00002615",
X"00003360",
X"0000262a",
X"00003351",
X"0000263e",
X"00003341",
X"00002652",
X"00003332",
X"00002666",
X"00003323",
X"0000267a",
X"00003314",
X"0000268e",
X"00003304",
X"000026a2",
X"000032f5",
X"000026b6",
X"000032e6",
X"000026ca",
X"000032d7",
X"000026de",
X"000032c7",
X"000026f2",
X"000032b8",
X"00002706",
X"000032a9",
X"0000271a",
X"0000329a",
X"0000272e",
X"0000328a",
X"00002742",
X"0000327b",
X"00002756",
X"0000326c",
X"00002769",
X"0000325c",
X"0000277d",
X"0000324c",
X"00002791",
X"0000323d",
X"000027a4",
X"0000322d",
X"000027b8",
X"0000321d",
X"000027cb",
X"0000320e",
X"000027df",
X"000031fe",
X"000027f3",
X"000031ee",
X"00002806",
X"000031de",
X"0000281a",
X"000031cf",
X"0000282e",
X"000031bf",
X"00002841",
X"000031af",
X"00002855",
X"000031a0",
X"00002868",
X"00003190",
X"0000287c",
X"00003180",
X"00002890",
X"00003170",
X"000028a3",
X"00003160",
X"000028b6",
X"00003150",
X"000028ca",
X"00003140",
X"000028dd",
X"00003130",
X"000028f0",
X"0000311f",
X"00002903",
X"0000310f",
X"00002917",
X"000030ff",
X"0000292a",
X"000030ef",
X"0000293d",
X"000030df",
X"00002950",
X"000030cf",
X"00002964",
X"000030be",
X"00002977",
X"000030ae",
X"0000298a",
X"0000309e",
X"0000299d",
X"0000308e",
X"000029b1",
X"0000307e",
X"000029c4",
X"0000306d",
X"000029d7",
X"0000305d",
X"000029ea",
X"0000304c",
X"000029fd",
X"0000303b",
X"00002a0f",
X"0000302b",
X"00002a22",
X"0000301a",
X"00002a35",
X"00003009",
X"00002a48",
X"00002ff9",
X"00002a5b",
X"00002fe8",
X"00002a6d",
X"00002fd8",
X"00002a80",
X"00002fc7",
X"00002a93",
X"00002fb6",
X"00002aa6",
X"00002fa6",
X"00002ab9",
X"00002f95",
X"00002acb",
X"00002f84",
X"00002ade",
X"00002f74",
X"00002af1",
X"00002f63",
X"00002b04",
X"00002f52",
X"00002b16",
X"00002f41",
X"00002b28",
X"00002f30",
X"00002b3b",
X"00002f1e",
X"00002b4d",
X"00002f0d",
X"00002b60",
X"00002efc",
X"00002b72",
X"00002eeb",
X"00002b84",
X"00002eda",
X"00002b97",
X"00002ec9",
X"00002ba9",
X"00002eb8",
X"00002bbb",
X"00002ea7",
X"00002bce",
X"00002e95",
X"00002be0",
X"00002e84",
X"00002bf3",
X"00002e73",
X"00002c05",
X"00002e62",
X"00002c17",
X"00002e51",
X"00002c2a",
X"00002e3f",
X"00002c3c",
X"00002e2e",
X"00002c4e",
X"00002e1c",
X"00002c60",
X"00002e0a",
X"00002c72",
X"00002df9",
X"00002c84",
X"00002de7",
X"00002c96",
X"00002dd6",
X"00002ca8",
X"00002dc4",
X"00002cba",
X"00002db3",
X"00002ccc",
X"00002da1",
X"00002cde",
X"00002d90",
X"00002cf0",
X"00002d7e",
X"00002d02",
X"00002d6c",
X"00002d14",
X"00002d5b",
X"00002d26",
X"00002d49",
X"00002d38",
X"00001fff",
X"ffffffe7",
X"00001fff",
X"ffffffb5",
X"00001ffe",
X"ffffff83",
X"00001ffd",
X"ffffff51",
X"00001ffc",
X"ffffff1e",
X"00001ffa",
X"fffffeec",
X"00001ff8",
X"fffffeba",
X"00001ff6",
X"fffffe88",
X"00001ff4",
X"fffffe55",
X"00001ff1",
X"fffffe23",
X"00001fee",
X"fffffdf1",
X"00001feb",
X"fffffdbf",
X"00001fe7",
X"fffffd8d",
X"00001fe3",
X"fffffd5b",
X"00001fdf",
X"fffffd29",
X"00001fda",
X"fffffcf7",
X"00001fd5",
X"fffffcc4",
X"00001fd0",
X"fffffc92",
X"00001fca",
X"fffffc60",
X"00001fc5",
X"fffffc2e",
X"00001fbf",
X"fffffbfd",
X"00001fb8",
X"fffffbcb",
X"00001fb1",
X"fffffb99",
X"00001faa",
X"fffffb67",
X"00001fa3",
X"fffffb36",
X"00001f9b",
X"fffffb04",
X"00001f93",
X"fffffad2",
X"00001f8b",
X"fffffaa1",
X"00001f82",
X"fffffa6f",
X"00001f79",
X"fffffa3e",
X"00001f70",
X"fffffa0d",
X"00001f67",
X"fffff9db",
X"00001f5d",
X"fffff9aa",
X"00001f52",
X"fffff979",
X"00001f48",
X"fffff947",
X"00001f3e",
X"fffff916",
X"00001f33",
X"fffff8e5",
X"00001f27",
X"fffff8b4",
X"00001f1b",
X"fffff883",
X"00001f10",
X"fffff852",
X"00001f04",
X"fffff822",
X"00001ef7",
X"fffff7f1",
X"00001eea",
X"fffff7c0",
X"00001edd",
X"fffff790",
X"00001ed0",
X"fffff75f",
X"00001ec2",
X"fffff72f",
X"00001eb4",
X"fffff6ff",
X"00001ea6",
X"fffff6cf",
X"00001e97",
X"fffff69f",
X"00001e88",
X"fffff66f",
X"00001e79",
X"fffff63f",
X"00001e6a",
X"fffff60f",
X"00001e5a",
X"fffff5df",
X"00001e49",
X"fffff5b0",
X"00001e39",
X"fffff580",
X"00001e29",
X"fffff550",
X"00001e18",
X"fffff521",
X"00001e06",
X"fffff4f2",
X"00001df5",
X"fffff4c3",
X"00001de3",
X"fffff494",
X"00001dd1",
X"fffff465",
X"00001dbf",
X"fffff436",
X"00001dac",
X"fffff407",
X"00001d99",
X"fffff3d9",
X"00001d86",
X"fffff3aa",
X"00001d72",
X"fffff37c",
X"00001d5e",
X"fffff34e",
X"00001d4a",
X"fffff320",
X"00001d36",
X"fffff2f2",
X"00001d21",
X"fffff2c4",
X"00001d0c",
X"fffff297",
X"00001cf7",
X"fffff269",
X"00001ce2",
X"fffff23b",
X"00001ccc",
X"fffff20e",
X"00001cb6",
X"fffff1e1",
X"00001ca0",
X"fffff1b4",
X"00001c89",
X"fffff187",
X"00001c72",
X"fffff15b",
X"00001c5b",
X"fffff12e",
X"00001c44",
X"fffff101",
X"00001c2c",
X"fffff0d5",
X"00001c14",
X"fffff0a9",
X"00001bfc",
X"fffff07d",
X"00001be4",
X"fffff051",
X"00001bcb",
X"fffff025",
X"00001bb1",
X"ffffeff9",
X"00001b98",
X"ffffefce",
X"00001b7f",
X"ffffefa3",
X"00001b65",
X"ffffef78",
X"00001b4a",
X"ffffef4d",
X"00001b30",
X"ffffef22",
X"00001b16",
X"ffffeef7",
X"00001afb",
X"ffffeecd",
X"00001adf",
X"ffffeea3",
X"00001ac4",
X"ffffee79",
X"00001aa9",
X"ffffee4f",
X"00001a8d",
X"ffffee25",
X"00001a70",
X"ffffedfb",
X"00001a54",
X"ffffedd2",
X"00001a37",
X"ffffeda8",
X"00001a1a",
X"ffffed7f",
X"000019fd",
X"ffffed56",
X"000019e0",
X"ffffed2e",
X"000019c2",
X"ffffed05",
X"000019a4",
X"ffffecdc",
X"00001986",
X"ffffecb4",
X"00001967",
X"ffffec8c",
X"00001949",
X"ffffec64",
X"0000192a",
X"ffffec3d",
X"0000190a",
X"ffffec16",
X"000018eb",
X"ffffebee",
X"000018cc",
X"ffffebc7",
X"000018ac",
X"ffffeba0",
X"0000188b",
X"ffffeb7a",
X"0000186b",
X"ffffeb53",
X"0000184b",
X"ffffeb2d",
X"0000182a",
X"ffffeb07",
X"00001809",
X"ffffeae1",
X"000017e7",
X"ffffeabb",
X"000017c6",
X"ffffea96",
X"000017a4",
X"ffffea71",
X"00001782",
X"ffffea4c",
X"00001760",
X"ffffea27",
X"0000173e",
X"ffffea02",
X"0000171b",
X"ffffe9de",
X"000016f8",
X"ffffe9ba",
X"000016d5",
X"ffffe996",
X"000016b2",
X"ffffe972",
X"0000168e",
X"ffffe94e",
X"0000166a",
X"ffffe92b",
X"00001646",
X"ffffe908",
X"00001622",
X"ffffe8e5",
X"000015fe",
X"ffffe8c2",
X"000015d9",
X"ffffe8a0",
X"000015b4",
X"ffffe87e",
X"0000158f",
X"ffffe85c",
X"0000156a",
X"ffffe83a",
X"00001545",
X"ffffe819",
X"0000151f",
X"ffffe7f7",
X"000014f9",
X"ffffe7d6",
X"000014d3",
X"ffffe7b5",
X"000014ad",
X"ffffe795",
X"00001486",
X"ffffe775",
X"00001460",
X"ffffe754",
X"00001439",
X"ffffe734",
X"00001412",
X"ffffe715",
X"000013ea",
X"ffffe6f6",
X"000013c3",
X"ffffe6d6",
X"0000139c",
X"ffffe6b7",
X"00001374",
X"ffffe699",
X"0000134c",
X"ffffe67a",
X"00001324",
X"ffffe65c",
X"000012fb",
X"ffffe63e",
X"000012d2",
X"ffffe620",
X"000012aa",
X"ffffe603",
X"00001281",
X"ffffe5e6",
X"00001258",
X"ffffe5c9",
X"0000122e",
X"ffffe5ac",
X"00001205",
X"ffffe590",
X"000011db",
X"ffffe573",
X"000011b1",
X"ffffe557",
X"00001187",
X"ffffe53c",
X"0000115d",
X"ffffe521",
X"00001133",
X"ffffe505",
X"00001109",
X"ffffe4ea",
X"000010de",
X"ffffe4d0",
X"000010b3",
X"ffffe4b6",
X"00001088",
X"ffffe49b",
X"0000105d",
X"ffffe481",
X"00001032",
X"ffffe468",
X"00001007",
X"ffffe44f",
X"00000fdb",
X"ffffe435",
X"00000faf",
X"ffffe41c",
X"00000f83",
X"ffffe404",
X"00000f57",
X"ffffe3ec",
X"00000f2b",
X"ffffe3d4",
X"00000eff",
X"ffffe3bc",
X"00000ed2",
X"ffffe3a5",
X"00000ea5",
X"ffffe38e",
X"00000e79",
X"ffffe377",
X"00000e4c",
X"ffffe360",
X"00000e1f",
X"ffffe34a",
X"00000df2",
X"ffffe334",
X"00000dc5",
X"ffffe31e",
X"00000d97",
X"ffffe309",
X"00000d69",
X"ffffe2f4",
X"00000d3c",
X"ffffe2df",
X"00000d0e",
X"ffffe2ca",
X"00000ce0",
X"ffffe2b6",
X"00000cb2",
X"ffffe2a2",
X"00000c84",
X"ffffe28e",
X"00000c56",
X"ffffe27a",
X"00000c27",
X"ffffe267",
X"00000bf9",
X"ffffe254",
X"00000bca",
X"ffffe241",
X"00000b9b",
X"ffffe22f",
X"00000b6c",
X"ffffe21d",
X"00000b3d",
X"ffffe20b",
X"00000b0e",
X"ffffe1fa",
X"00000adf",
X"ffffe1e8",
X"00000ab0",
X"ffffe1d7",
X"00000a80",
X"ffffe1c7",
X"00000a50",
X"ffffe1b7",
X"00000a21",
X"ffffe1a6",
X"000009f1",
X"ffffe196",
X"000009c1",
X"ffffe187",
X"00000991",
X"ffffe178",
X"00000961",
X"ffffe169",
X"00000931",
X"ffffe15a",
X"00000901",
X"ffffe14c",
X"000008d1",
X"ffffe13e",
X"000008a1",
X"ffffe130",
X"00000870",
X"ffffe123",
X"00000840",
X"ffffe116",
X"0000080f",
X"ffffe109",
X"000007de",
X"ffffe0fc",
X"000007ae",
X"ffffe0f0",
X"0000077d",
X"ffffe0e5",
X"0000074c",
X"ffffe0d9",
X"0000071b",
X"ffffe0cd",
X"000006ea",
X"ffffe0c2",
X"000006b9",
X"ffffe0b8",
X"00000687",
X"ffffe0ae",
X"00000656",
X"ffffe0a3",
X"00000625",
X"ffffe099",
X"000005f3",
X"ffffe090",
X"000005c2",
X"ffffe087",
X"00000591",
X"ffffe07e",
X"0000055f",
X"ffffe075",
X"0000052e",
X"ffffe06d",
X"000004fc",
X"ffffe065",
X"000004ca",
X"ffffe05d",
X"00000499",
X"ffffe056",
X"00000467",
X"ffffe04f",
X"00000435",
X"ffffe048",
X"00000403",
X"ffffe041",
X"000003d2",
X"ffffe03b",
X"000003a0",
X"ffffe036",
X"0000036e",
X"ffffe030",
X"0000033c",
X"ffffe02b",
X"00000309",
X"ffffe026",
X"000002d7",
X"ffffe021",
X"000002a5",
X"ffffe01d",
X"00000273",
X"ffffe019",
X"00000241",
X"ffffe015",
X"0000020f",
X"ffffe012",
X"000001dd",
X"ffffe00f",
X"000001ab",
X"ffffe00c",
X"00000178",
X"ffffe00a",
X"00000146",
X"ffffe008",
X"00000114",
X"ffffe006",
X"000000e2",
X"ffffe004",
X"000000af",
X"ffffe003",
X"0000007d",
X"ffffe002",
X"0000004b",
X"ffffe001",
X"00000019",
X"ffffe001"
);
end;


