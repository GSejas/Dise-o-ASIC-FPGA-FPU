n = 256

bitrev:
0: "126"
1: "0"
2: "62"
3: "64"
4: "94"
5: "32"
6: "30"
7: "96"
8: "110"
9: "16"
10: "46"
11: "80"
12: "78"
13: "48"
14: "14"
15: "112"
16: "118"
17: "8"
18: "54"
19: "72"
20: "86"
21: "40"
22: "22"
23: "104"
24: "102"
25: "24"
26: "38"
27: "88"
28: "70"
29: "56"
30: "6"
31: "120"
32: "122"
33: "4"
34: "58"
35: "68"
36: "90"
37: "36"
38: "26"
39: "100"
40: "106"
41: "20"
42: "42"
43: "84"
44: "74"
45: "52"
46: "10"
47: "116"
48: "114"
49: "12"
50: "50"
51: "76"
52: "82"
53: "44"
54: "18"
55: "108"
56: "98"
57: "28"
58: "34"
59: "92"
60: "66"
61: "60"
62: "2"
63: "124"
T:
X"4000", 
X"0", 
X"3fec", 
X"fffffcdc", 
X"3fb1", 
X"fffff9ba", 
X"3f4f", 
X"fffff69c", 
X"3ec5", 
X"fffff384", 
X"3e15", 
X"fffff073", 
X"3d3f", 
X"ffffed6c", 
X"3c42", 
X"ffffea70", 
X"3b21", 
X"ffffe782", 
X"39db", 
X"ffffe4a3", 
X"3871", 
X"ffffe1d5", 
X"36e5", 
X"ffffdf19", 
X"3537", 
X"ffffdc72", 
X"3368", 
X"ffffd9e0", 
X"3179", 
X"ffffd766", 
X"2f6c", 
X"ffffd505", 
X"2d41", 
X"ffffd2bf", 
X"2afb", 
X"ffffd094", 
X"289a", 
X"ffffce87", 
X"2620", 
X"ffffcc98", 
X"238e", 
X"ffffcac9", 
X"20e7", 
X"ffffc91b", 
X"1e2b", 
X"ffffc78f", 
X"1b5d", 
X"ffffc625", 
X"187e", 
X"ffffc4df", 
X"1590", 
X"ffffc3be", 
X"1294", 
X"ffffc2c1", 
X"f8d", 
X"ffffc1eb", 
X"c7c", 
X"ffffc13b", 
X"964", 
X"ffffc0b1", 
X"646", 
X"ffffc04f", 
X"324", 
X"ffffc014", 
X"0", 
X"ffffc000", 
X"fffffcdd", 
X"ffffc014", 
X"fffff9bb", 
X"ffffc04f", 
X"fffff69d", 
X"ffffc0b1", 
X"fffff385", 
X"ffffc13b", 
X"fffff074", 
X"ffffc1eb", 
X"ffffed6d", 
X"ffffc2c1", 
X"ffffea71", 
X"ffffc3be", 
X"ffffe783", 
X"ffffc4df", 
X"ffffe4a4", 
X"ffffc625", 
X"ffffe1d6", 
X"ffffc78f", 
X"ffffdf1a", 
X"ffffc91b", 
X"ffffdc73", 
X"ffffcac9", 
X"ffffd9e1", 
X"ffffcc98", 
X"ffffd767", 
X"ffffce87", 
X"ffffd506", 
X"ffffd094", 
X"ffffd2c0", 
X"ffffd2bf", 
X"ffffd095", 
X"ffffd505", 
X"ffffce88", 
X"ffffd766", 
X"ffffcc99", 
X"ffffd9e0", 
X"ffffcaca", 
X"ffffdc72", 
X"ffffc91c", 
X"ffffdf19", 
X"ffffc790", 
X"ffffe1d5", 
X"ffffc626", 
X"ffffe4a3", 
X"ffffc4e0", 
X"ffffe782", 
X"ffffc3bf", 
X"ffffea70", 
X"ffffc2c2", 
X"ffffed6c", 
X"ffffc1ec", 
X"fffff073", 
X"ffffc13c", 
X"fffff384", 
X"ffffc0b2", 
X"fffff69c", 
X"ffffc050", 
X"fffff9ba", 
X"ffffc015", 
X"fffffcdc", 
X"3ffe", 
X"64", 
X"3ffc", 
X"12d", 
X"3ff7", 
X"1f6", 
X"3fef", 
X"2bf", 
X"3fe6", 
X"388", 
X"3fda", 
X"450", 
X"3fcb", 
X"519", 
X"3fb9", 
X"5e1", 
X"3fa6", 
X"6aa", 
X"3f90", 
X"772", 
X"3f77", 
X"839", 
X"3f5c", 
X"900", 
X"3f3f", 
X"9c7", 
X"3f1f", 
X"a8d", 
X"3efc", 
X"b53", 
X"3ed7", 
X"c19", 
X"3eb0", 
X"cde", 
X"3e86", 
X"da3", 
X"3e5a", 
X"e67", 
X"3e2c", 
X"f2b", 
X"3dfb", 
X"fee", 
X"3dc8", 
X"10b0", 
X"3d93", 
X"1172", 
X"3d5b", 
X"1233", 
X"3d20", 
X"12f3", 
X"3ce3", 
X"13b3", 
X"3ca4", 
X"1472", 
X"3c62", 
X"1530", 
X"3c1f", 
X"15ee", 
X"3bd9", 
X"16aa", 
X"3b90", 
X"1766", 
X"3b46", 
X"1820", 
X"3af9", 
X"18da", 
X"3aa9", 
X"1992", 
X"3a58", 
X"1a4a", 
X"3a04", 
X"1b01", 
X"39af", 
X"1bb7", 
X"3957", 
X"1c6b", 
X"38fc", 
X"1d1f", 
X"389f", 
X"1dd1", 
X"3840", 
X"1e83", 
X"37e0", 
X"1f33", 
X"377d", 
X"1fe2", 
X"3717", 
X"2090", 
X"36b0", 
X"213c", 
X"3646", 
X"21e7", 
X"35db", 
X"2291", 
X"356d", 
X"2339", 
X"34fe", 
X"23e1", 
X"348c", 
X"2487", 
X"3418", 
X"252b", 
X"33a2", 
X"25ce", 
X"332b", 
X"2670", 
X"32b1", 
X"2710", 
X"3235", 
X"27ae", 
X"31b7", 
X"284b", 
X"3138", 
X"28e7", 
X"30b6", 
X"2981", 
X"3033", 
X"2a19", 
X"2fae", 
X"2aaf", 
X"2f27", 
X"2b44", 
X"2e9e", 
X"2bd7", 
X"2e13", 
X"2c69", 
X"2d87", 
X"2cf9", 
X"1ffd", 
X"ffffff37", 
X"1fea", 
X"fffffda6", 
X"1fc2", 
X"fffffc15", 
X"1f87", 
X"fffffa88", 
X"1f39", 
X"fffff8fd", 
X"1ed7", 
X"fffff777", 
X"1e62", 
X"fffff5f7", 
X"1ddb", 
X"fffff47c", 
X"1d41", 
X"fffff309", 
X"1c95", 
X"fffff19d", 
X"1bd8", 
X"fffff03a", 
X"1b09", 
X"ffffeee2", 
X"1a29", 
X"ffffed93", 
X"193a", 
X"ffffec50", 
X"183b", 
X"ffffeb19", 
X"172d", 
X"ffffe9f0", 
X"1610", 
X"ffffe8d3", 
X"14e7", 
X"ffffe7c5", 
X"13b0", 
X"ffffe6c6", 
X"126d", 
X"ffffe5d7", 
X"111e", 
X"ffffe4f7", 
X"fc6", 
X"ffffe428", 
X"e63", 
X"ffffe36b", 
X"cf7", 
X"ffffe2bf", 
X"b84", 
X"ffffe225", 
X"a09", 
X"ffffe19e", 
X"889", 
X"ffffe129", 
X"703", 
X"ffffe0c7", 
X"578", 
X"ffffe079", 
X"3eb", 
X"ffffe03e", 
X"25a", 
X"ffffe016", 
X"c9", 
X"ffffe003", 

