`ifndef __XC3S_RAM16X233_D_V__
`define __XC3S_RAM16X233_D_V__

//`include "RAM16X1D.v"

module XC3S_RAM16X233_D (DIN, ADDR1, ADDR2, WE, WCLK, O_DOUT1, O_DOUT2);

parameter data_width = 233;//Replace with desired data-bus width 
                         
input wire [232:0]DIN;
input wire [3:0] ADDR1, ADDR2;
input wire WE;
input wire WCLK;

output wire [232:0]O_DOUT1, O_DOUT2;

wire [232:0]DOUT1, DOUT2;


/*Remember to Instantiate a Distributed SelectRAM block for each Data port
  and to give each instance a unique name...The following is an example of instantiation 
  for a 16 X 8-bit RAM. */
RAM16X1D U_RAM16X1D_0(DOUT2[0], DOUT1[0], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[0], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_1(DOUT2[1], DOUT1[1], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[1], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_2(DOUT2[2], DOUT1[2], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[2], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_3(DOUT2[3], DOUT1[3], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[3], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_4(DOUT2[4], DOUT1[4], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[4], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_5(DOUT2[5], DOUT1[5], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[5], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_6(DOUT2[6], DOUT1[6], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[6], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_7(DOUT2[7], DOUT1[7], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[7], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_8(DOUT2[8], DOUT1[8], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[8], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_9(DOUT2[9], DOUT1[9], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[9], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);

RAM16X1D U_RAM16X1D_10(DOUT2[10], DOUT1[10], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[10], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_11(DOUT2[11], DOUT1[11], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[11], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_12(DOUT2[12], DOUT1[12], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[12], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_13(DOUT2[13], DOUT1[13], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[13], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_14(DOUT2[14], DOUT1[14], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[14], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_15(DOUT2[15], DOUT1[15], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[15], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_16(DOUT2[16], DOUT1[16], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[16], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_17(DOUT2[17], DOUT1[17], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[17], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_18(DOUT2[18], DOUT1[18], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[18], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_19(DOUT2[19], DOUT1[19], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[19], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);

RAM16X1D U_RAM16X1D_20(DOUT2[20], DOUT1[20], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[20], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_21(DOUT2[21], DOUT1[21], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[21], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_22(DOUT2[22], DOUT1[22], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[22], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_23(DOUT2[23], DOUT1[23], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[23], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_24(DOUT2[24], DOUT1[24], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[24], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_25(DOUT2[25], DOUT1[25], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[25], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_26(DOUT2[26], DOUT1[26], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[26], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_27(DOUT2[27], DOUT1[27], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[27], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_28(DOUT2[28], DOUT1[28], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[28], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_29(DOUT2[29], DOUT1[29], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[29], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);

RAM16X1D U_RAM16X1D_30(DOUT2[30], DOUT1[30], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[30], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_31(DOUT2[31], DOUT1[31], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[31], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_32(DOUT2[32], DOUT1[32], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[32], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_33(DOUT2[33], DOUT1[33], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[33], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_34(DOUT2[34], DOUT1[34], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[34], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_35(DOUT2[35], DOUT1[35], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[35], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_36(DOUT2[36], DOUT1[36], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[36], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_37(DOUT2[37], DOUT1[37], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[37], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_38(DOUT2[38], DOUT1[38], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[38], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_39(DOUT2[39], DOUT1[39], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[39], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);

RAM16X1D U_RAM16X1D_40(DOUT2[40], DOUT1[40], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[40], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_41(DOUT2[41], DOUT1[41], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[41], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_42(DOUT2[42], DOUT1[42], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[42], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_43(DOUT2[43], DOUT1[43], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[43], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_44(DOUT2[44], DOUT1[44], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[44], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_45(DOUT2[45], DOUT1[45], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[45], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_46(DOUT2[46], DOUT1[46], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[46], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_47(DOUT2[47], DOUT1[47], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[47], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_48(DOUT2[48], DOUT1[48], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[48], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_49(DOUT2[49], DOUT1[49], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[49], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);

RAM16X1D U_RAM16X1D_50(DOUT2[50], DOUT1[50], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[50], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_51(DOUT2[51], DOUT1[51], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[51], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_52(DOUT2[52], DOUT1[52], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[52], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_53(DOUT2[53], DOUT1[53], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[53], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_54(DOUT2[54], DOUT1[54], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[54], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_55(DOUT2[55], DOUT1[55], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[55], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_56(DOUT2[56], DOUT1[56], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[56], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_57(DOUT2[57], DOUT1[57], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[57], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_58(DOUT2[58], DOUT1[58], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[58], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_59(DOUT2[59], DOUT1[59], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[59], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);

RAM16X1D U_RAM16X1D_60(DOUT2[60], DOUT1[60], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[60], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_61(DOUT2[61], DOUT1[61], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[61], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_62(DOUT2[62], DOUT1[62], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[62], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_63(DOUT2[63], DOUT1[63], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[63], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_64(DOUT2[64], DOUT1[64], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[64], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_65(DOUT2[65], DOUT1[65], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[65], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_66(DOUT2[66], DOUT1[66], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[66], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_67(DOUT2[67], DOUT1[67], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[67], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_68(DOUT2[68], DOUT1[68], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[68], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_69(DOUT2[69], DOUT1[69], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[69], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);

RAM16X1D U_RAM16X1D_70(DOUT2[70], DOUT1[70], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[70], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_71(DOUT2[71], DOUT1[71], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[71], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_72(DOUT2[72], DOUT1[72], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[72], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_73(DOUT2[73], DOUT1[73], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[73], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_74(DOUT2[74], DOUT1[74], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[74], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_75(DOUT2[75], DOUT1[75], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[75], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_76(DOUT2[76], DOUT1[76], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[76], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_77(DOUT2[77], DOUT1[77], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[77], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_78(DOUT2[78], DOUT1[78], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[78], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_79(DOUT2[79], DOUT1[79], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[79], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);

RAM16X1D U_RAM16X1D_80(DOUT2[80], DOUT1[80], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[80], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_81(DOUT2[81], DOUT1[81], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[81], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_82(DOUT2[82], DOUT1[82], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[82], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_83(DOUT2[83], DOUT1[83], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[83], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_84(DOUT2[84], DOUT1[84], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[84], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_85(DOUT2[85], DOUT1[85], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[85], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_86(DOUT2[86], DOUT1[86], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[86], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_87(DOUT2[87], DOUT1[87], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[87], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_88(DOUT2[88], DOUT1[88], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[88], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_89(DOUT2[89], DOUT1[89], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[89], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);

RAM16X1D U_RAM16X1D_90(DOUT2[90], DOUT1[90], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[90], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_91(DOUT2[91], DOUT1[91], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[91], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_92(DOUT2[92], DOUT1[92], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[92], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_93(DOUT2[93], DOUT1[93], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[93], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_94(DOUT2[94], DOUT1[94], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[94], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_95(DOUT2[95], DOUT1[95], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[95], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_96(DOUT2[96], DOUT1[96], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[96], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_97(DOUT2[97], DOUT1[97], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[97], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_98(DOUT2[98], DOUT1[98], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[98], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_99(DOUT2[99], DOUT1[99], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[99], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);

RAM16X1D U_RAM16X1D_100(DOUT2[100], DOUT1[100], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[100], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_101(DOUT2[101], DOUT1[101], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[101], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_102(DOUT2[102], DOUT1[102], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[102], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_103(DOUT2[103], DOUT1[103], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[103], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_104(DOUT2[104], DOUT1[104], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[104], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_105(DOUT2[105], DOUT1[105], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[105], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_106(DOUT2[106], DOUT1[106], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[106], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_107(DOUT2[107], DOUT1[107], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[107], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_108(DOUT2[108], DOUT1[108], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[108], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_109(DOUT2[109], DOUT1[109], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[109], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);

RAM16X1D U_RAM16X1D_110(DOUT2[110], DOUT1[110], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[110], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_111(DOUT2[111], DOUT1[111], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[111], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_112(DOUT2[112], DOUT1[112], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[112], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_113(DOUT2[113], DOUT1[113], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[113], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_114(DOUT2[114], DOUT1[114], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[114], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_115(DOUT2[115], DOUT1[115], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[115], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_116(DOUT2[116], DOUT1[116], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[116], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_117(DOUT2[117], DOUT1[117], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[117], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_118(DOUT2[118], DOUT1[118], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[118], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_119(DOUT2[119], DOUT1[119], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[119], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);

RAM16X1D U_RAM16X1D_120(DOUT2[120], DOUT1[120], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[120], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_121(DOUT2[121], DOUT1[121], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[121], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_122(DOUT2[122], DOUT1[122], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[122], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_123(DOUT2[123], DOUT1[123], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[123], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_124(DOUT2[124], DOUT1[124], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[124], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_125(DOUT2[125], DOUT1[125], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[125], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_126(DOUT2[126], DOUT1[126], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[126], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_127(DOUT2[127], DOUT1[127], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[127], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_128(DOUT2[128], DOUT1[128], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[128], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_129(DOUT2[129], DOUT1[129], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[129], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);

RAM16X1D U_RAM16X1D_130(DOUT2[130], DOUT1[130], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[130], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_131(DOUT2[131], DOUT1[131], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[131], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_132(DOUT2[132], DOUT1[132], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[132], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_133(DOUT2[133], DOUT1[133], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[133], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_134(DOUT2[134], DOUT1[134], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[134], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_135(DOUT2[135], DOUT1[135], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[135], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_136(DOUT2[136], DOUT1[136], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[136], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_137(DOUT2[137], DOUT1[137], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[137], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_138(DOUT2[138], DOUT1[138], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[138], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_139(DOUT2[139], DOUT1[139], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[139], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);

RAM16X1D U_RAM16X1D_140(DOUT2[140], DOUT1[140], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[140], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_141(DOUT2[141], DOUT1[141], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[141], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_142(DOUT2[142], DOUT1[142], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[142], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_143(DOUT2[143], DOUT1[143], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[143], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_144(DOUT2[144], DOUT1[144], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[144], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_145(DOUT2[145], DOUT1[145], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[145], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_146(DOUT2[146], DOUT1[146], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[146], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_147(DOUT2[147], DOUT1[147], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[147], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_148(DOUT2[148], DOUT1[148], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[148], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_149(DOUT2[149], DOUT1[149], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[149], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);

RAM16X1D U_RAM16X1D_150(DOUT2[150], DOUT1[150], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[150], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_151(DOUT2[151], DOUT1[151], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[151], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_152(DOUT2[152], DOUT1[152], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[152], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_153(DOUT2[153], DOUT1[153], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[153], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_154(DOUT2[154], DOUT1[154], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[154], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_155(DOUT2[155], DOUT1[155], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[155], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_156(DOUT2[156], DOUT1[156], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[156], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_157(DOUT2[157], DOUT1[157], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[157], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_158(DOUT2[158], DOUT1[158], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[158], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_159(DOUT2[159], DOUT1[159], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[159], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);

RAM16X1D U_RAM16X1D_160(DOUT2[160], DOUT1[160], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[160], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_161(DOUT2[161], DOUT1[161], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[161], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_162(DOUT2[162], DOUT1[162], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[162], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_163(DOUT2[163], DOUT1[163], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[163], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_164(DOUT2[164], DOUT1[164], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[164], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_165(DOUT2[165], DOUT1[165], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[165], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_166(DOUT2[166], DOUT1[166], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[166], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_167(DOUT2[167], DOUT1[167], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[167], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_168(DOUT2[168], DOUT1[168], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[168], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_169(DOUT2[169], DOUT1[169], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[169], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);

RAM16X1D U_RAM16X1D_170(DOUT2[170], DOUT1[170], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[170], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_171(DOUT2[171], DOUT1[171], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[171], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_172(DOUT2[172], DOUT1[172], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[172], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_173(DOUT2[173], DOUT1[173], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[173], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_174(DOUT2[174], DOUT1[174], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[174], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_175(DOUT2[175], DOUT1[175], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[175], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_176(DOUT2[176], DOUT1[176], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[176], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_177(DOUT2[177], DOUT1[177], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[177], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_178(DOUT2[178], DOUT1[178], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[178], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_179(DOUT2[179], DOUT1[179], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[179], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);

RAM16X1D U_RAM16X1D_180(DOUT2[180], DOUT1[180], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[180], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_181(DOUT2[181], DOUT1[181], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[181], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_182(DOUT2[182], DOUT1[182], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[182], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_183(DOUT2[183], DOUT1[183], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[183], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_184(DOUT2[184], DOUT1[184], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[184], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_185(DOUT2[185], DOUT1[185], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[185], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_186(DOUT2[186], DOUT1[186], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[186], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_187(DOUT2[187], DOUT1[187], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[187], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_188(DOUT2[188], DOUT1[188], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[188], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_189(DOUT2[189], DOUT1[189], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[189], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);

RAM16X1D U_RAM16X1D_190(DOUT2[190], DOUT1[190], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[190], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_191(DOUT2[191], DOUT1[191], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[191], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_192(DOUT2[192], DOUT1[192], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[192], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_193(DOUT2[193], DOUT1[193], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[193], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_194(DOUT2[194], DOUT1[194], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[194], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_195(DOUT2[195], DOUT1[195], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[195], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_196(DOUT2[196], DOUT1[196], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[196], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_197(DOUT2[197], DOUT1[197], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[197], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_198(DOUT2[198], DOUT1[198], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[198], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_199(DOUT2[199], DOUT1[199], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[199], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);

RAM16X1D U_RAM16X1D_200(DOUT2[200], DOUT1[200], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[200], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_201(DOUT2[201], DOUT1[201], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[201], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_202(DOUT2[202], DOUT1[202], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[202], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_203(DOUT2[203], DOUT1[203], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[203], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_204(DOUT2[204], DOUT1[204], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[204], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_205(DOUT2[205], DOUT1[205], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[205], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_206(DOUT2[206], DOUT1[206], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[206], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_207(DOUT2[207], DOUT1[207], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[207], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_208(DOUT2[208], DOUT1[208], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[208], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_209(DOUT2[209], DOUT1[209], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[209], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);

RAM16X1D U_RAM16X1D_210(DOUT2[210], DOUT1[210], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[210], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_211(DOUT2[211], DOUT1[211], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[211], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_212(DOUT2[212], DOUT1[212], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[212], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_213(DOUT2[213], DOUT1[213], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[213], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_214(DOUT2[214], DOUT1[214], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[214], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_215(DOUT2[215], DOUT1[215], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[215], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_216(DOUT2[216], DOUT1[216], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[216], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_217(DOUT2[217], DOUT1[217], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[217], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_218(DOUT2[218], DOUT1[218], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[218], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_219(DOUT2[219], DOUT1[219], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[219], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);

RAM16X1D U_RAM16X1D_220(DOUT2[220], DOUT1[220], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[220], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_221(DOUT2[221], DOUT1[221], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[221], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_222(DOUT2[222], DOUT1[222], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[222], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_223(DOUT2[223], DOUT1[223], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[223], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_224(DOUT2[224], DOUT1[224], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[224], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_225(DOUT2[225], DOUT1[225], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[225], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_226(DOUT2[226], DOUT1[226], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[226], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_227(DOUT2[227], DOUT1[227], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[227], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_228(DOUT2[228], DOUT1[228], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[228], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_229(DOUT2[229], DOUT1[229], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[229], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);

RAM16X1D U_RAM16X1D_230(DOUT2[230], DOUT1[230], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[230], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_231(DOUT2[231], DOUT1[231], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[231], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);
RAM16X1D U_RAM16X1D_232(DOUT2[232], DOUT1[232], ADDR1[0], ADDR1[1], ADDR1[2], ADDR1[3], DIN[232], ADDR2[0], ADDR2[1], ADDR2[2], ADDR2[3], WCLK, WE);

//always @(posedge WCLK)
//begin
assign  O_DOUT1 = DOUT1;
assign  O_DOUT2 = DOUT2;
//end
endmodule

`endif
