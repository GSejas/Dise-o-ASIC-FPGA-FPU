/*******************************************************
* File Name     : hdl/ks26.v
* Module Name   : Karatsuba Multiplier
* Author        : Chester Rebeiro
* Institute     : Indian Institute of Technology, Madras
* Creation Time : 

* Comment       : Automatically generated from general.c
********************************************************/
`ifndef __KS_26_V__
`define __KS_26_V__

module ks26(a, b, d);

input wire [0:25] a;
input wire [0:25] b;
output wire [0:50] d;

wire m0, m1, m2, m3, m4, m5, m6, m7, m8, m9, m10, m11, m12, m13, m14, m15, m16, m17, m18, m19, m20, m21, m22, m23, m24, m25;
wire m0_1, m0_2, m0_3, m0_4, m0_5, m0_6, m0_7, m0_8, m0_9, m0_10, m0_11, m0_12, m0_13, m0_14, m0_15, m0_16, m0_17, m0_18, m0_19, m0_20, m0_21, m0_22, m0_23, m0_24, m0_25;
wire m1_2, m1_3, m1_4, m1_5, m1_6, m1_7, m1_8, m1_9, m1_10, m1_11, m1_12, m1_13, m1_14, m1_15, m1_16, m1_17, m1_18, m1_19, m1_20, m1_21, m1_22, m1_23, m1_24, m1_25;
wire m2_3, m2_4, m2_5, m2_6, m2_7, m2_8, m2_9, m2_10, m2_11, m2_12, m2_13, m2_14, m2_15, m2_16, m2_17, m2_18, m2_19, m2_20, m2_21, m2_22, m2_23, m2_24, m2_25;
wire m3_4, m3_5, m3_6, m3_7, m3_8, m3_9, m3_10, m3_11, m3_12, m3_13, m3_14, m3_15, m3_16, m3_17, m3_18, m3_19, m3_20, m3_21, m3_22, m3_23, m3_24, m3_25;
wire m4_5, m4_6, m4_7, m4_8, m4_9, m4_10, m4_11, m4_12, m4_13, m4_14, m4_15, m4_16, m4_17, m4_18, m4_19, m4_20, m4_21, m4_22, m4_23, m4_24, m4_25;
wire m5_6, m5_7, m5_8, m5_9, m5_10, m5_11, m5_12, m5_13, m5_14, m5_15, m5_16, m5_17, m5_18, m5_19, m5_20, m5_21, m5_22, m5_23, m5_24, m5_25;
wire m6_7, m6_8, m6_9, m6_10, m6_11, m6_12, m6_13, m6_14, m6_15, m6_16, m6_17, m6_18, m6_19, m6_20, m6_21, m6_22, m6_23, m6_24, m6_25;
wire m7_8, m7_9, m7_10, m7_11, m7_12, m7_13, m7_14, m7_15, m7_16, m7_17, m7_18, m7_19, m7_20, m7_21, m7_22, m7_23, m7_24, m7_25;
wire m8_9, m8_10, m8_11, m8_12, m8_13, m8_14, m8_15, m8_16, m8_17, m8_18, m8_19, m8_20, m8_21, m8_22, m8_23, m8_24, m8_25;
wire m9_10, m9_11, m9_12, m9_13, m9_14, m9_15, m9_16, m9_17, m9_18, m9_19, m9_20, m9_21, m9_22, m9_23, m9_24, m9_25;
wire m10_11, m10_12, m10_13, m10_14, m10_15, m10_16, m10_17, m10_18, m10_19, m10_20, m10_21, m10_22, m10_23, m10_24, m10_25;
wire m11_12, m11_13, m11_14, m11_15, m11_16, m11_17, m11_18, m11_19, m11_20, m11_21, m11_22, m11_23, m11_24, m11_25;
wire m12_13, m12_14, m12_15, m12_16, m12_17, m12_18, m12_19, m12_20, m12_21, m12_22, m12_23, m12_24, m12_25;
wire m13_14, m13_15, m13_16, m13_17, m13_18, m13_19, m13_20, m13_21, m13_22, m13_23, m13_24, m13_25;
wire m14_15, m14_16, m14_17, m14_18, m14_19, m14_20, m14_21, m14_22, m14_23, m14_24, m14_25;
wire m15_16, m15_17, m15_18, m15_19, m15_20, m15_21, m15_22, m15_23, m15_24, m15_25;
wire m16_17, m16_18, m16_19, m16_20, m16_21, m16_22, m16_23, m16_24, m16_25;
wire m17_18, m17_19, m17_20, m17_21, m17_22, m17_23, m17_24, m17_25;
wire m18_19, m18_20, m18_21, m18_22, m18_23, m18_24, m18_25;
wire m19_20, m19_21, m19_22, m19_23, m19_24, m19_25;
wire m20_21, m20_22, m20_23, m20_24, m20_25;
wire m21_22, m21_23, m21_24, m21_25;
wire m22_23, m22_24, m22_25;
wire m23_24, m23_25;
wire m24_25;
assign m0 = a[0] & b[0];
assign m1 = a[1] & b[1];
assign m2 = a[2] & b[2];
assign m3 = a[3] & b[3];
assign m4 = a[4] & b[4];
assign m5 = a[5] & b[5];
assign m6 = a[6] & b[6];
assign m7 = a[7] & b[7];
assign m8 = a[8] & b[8];
assign m9 = a[9] & b[9];
assign m10 = a[10] & b[10];
assign m11 = a[11] & b[11];
assign m12 = a[12] & b[12];
assign m13 = a[13] & b[13];
assign m14 = a[14] & b[14];
assign m15 = a[15] & b[15];
assign m16 = a[16] & b[16];
assign m17 = a[17] & b[17];
assign m18 = a[18] & b[18];
assign m19 = a[19] & b[19];
assign m20 = a[20] & b[20];
assign m21 = a[21] & b[21];
assign m22 = a[22] & b[22];
assign m23 = a[23] & b[23];
assign m24 = a[24] & b[24];
assign m25 = a[25] & b[25];
assign m0_1 = (a[0] ^ a[1]) & (b[0] ^ b[1]);
assign m0_2 = (a[0] ^ a[2]) & (b[0] ^ b[2]);
assign m0_3 = (a[0] ^ a[3]) & (b[0] ^ b[3]);
assign m0_4 = (a[0] ^ a[4]) & (b[0] ^ b[4]);
assign m0_5 = (a[0] ^ a[5]) & (b[0] ^ b[5]);
assign m0_6 = (a[0] ^ a[6]) & (b[0] ^ b[6]);
assign m0_7 = (a[0] ^ a[7]) & (b[0] ^ b[7]);
assign m0_8 = (a[0] ^ a[8]) & (b[0] ^ b[8]);
assign m0_9 = (a[0] ^ a[9]) & (b[0] ^ b[9]);
assign m0_10 = (a[0] ^ a[10]) & (b[0] ^ b[10]);
assign m0_11 = (a[0] ^ a[11]) & (b[0] ^ b[11]);
assign m0_12 = (a[0] ^ a[12]) & (b[0] ^ b[12]);
assign m0_13 = (a[0] ^ a[13]) & (b[0] ^ b[13]);
assign m0_14 = (a[0] ^ a[14]) & (b[0] ^ b[14]);
assign m0_15 = (a[0] ^ a[15]) & (b[0] ^ b[15]);
assign m0_16 = (a[0] ^ a[16]) & (b[0] ^ b[16]);
assign m0_17 = (a[0] ^ a[17]) & (b[0] ^ b[17]);
assign m0_18 = (a[0] ^ a[18]) & (b[0] ^ b[18]);
assign m0_19 = (a[0] ^ a[19]) & (b[0] ^ b[19]);
assign m0_20 = (a[0] ^ a[20]) & (b[0] ^ b[20]);
assign m0_21 = (a[0] ^ a[21]) & (b[0] ^ b[21]);
assign m0_22 = (a[0] ^ a[22]) & (b[0] ^ b[22]);
assign m0_23 = (a[0] ^ a[23]) & (b[0] ^ b[23]);
assign m0_24 = (a[0] ^ a[24]) & (b[0] ^ b[24]);
assign m0_25 = (a[0] ^ a[25]) & (b[0] ^ b[25]);
assign m1_2 = (a[1] ^ a[2]) & (b[1] ^ b[2]);
assign m1_3 = (a[1] ^ a[3]) & (b[1] ^ b[3]);
assign m1_4 = (a[1] ^ a[4]) & (b[1] ^ b[4]);
assign m1_5 = (a[1] ^ a[5]) & (b[1] ^ b[5]);
assign m1_6 = (a[1] ^ a[6]) & (b[1] ^ b[6]);
assign m1_7 = (a[1] ^ a[7]) & (b[1] ^ b[7]);
assign m1_8 = (a[1] ^ a[8]) & (b[1] ^ b[8]);
assign m1_9 = (a[1] ^ a[9]) & (b[1] ^ b[9]);
assign m1_10 = (a[1] ^ a[10]) & (b[1] ^ b[10]);
assign m1_11 = (a[1] ^ a[11]) & (b[1] ^ b[11]);
assign m1_12 = (a[1] ^ a[12]) & (b[1] ^ b[12]);
assign m1_13 = (a[1] ^ a[13]) & (b[1] ^ b[13]);
assign m1_14 = (a[1] ^ a[14]) & (b[1] ^ b[14]);
assign m1_15 = (a[1] ^ a[15]) & (b[1] ^ b[15]);
assign m1_16 = (a[1] ^ a[16]) & (b[1] ^ b[16]);
assign m1_17 = (a[1] ^ a[17]) & (b[1] ^ b[17]);
assign m1_18 = (a[1] ^ a[18]) & (b[1] ^ b[18]);
assign m1_19 = (a[1] ^ a[19]) & (b[1] ^ b[19]);
assign m1_20 = (a[1] ^ a[20]) & (b[1] ^ b[20]);
assign m1_21 = (a[1] ^ a[21]) & (b[1] ^ b[21]);
assign m1_22 = (a[1] ^ a[22]) & (b[1] ^ b[22]);
assign m1_23 = (a[1] ^ a[23]) & (b[1] ^ b[23]);
assign m1_24 = (a[1] ^ a[24]) & (b[1] ^ b[24]);
assign m1_25 = (a[1] ^ a[25]) & (b[1] ^ b[25]);
assign m2_3 = (a[2] ^ a[3]) & (b[2] ^ b[3]);
assign m2_4 = (a[2] ^ a[4]) & (b[2] ^ b[4]);
assign m2_5 = (a[2] ^ a[5]) & (b[2] ^ b[5]);
assign m2_6 = (a[2] ^ a[6]) & (b[2] ^ b[6]);
assign m2_7 = (a[2] ^ a[7]) & (b[2] ^ b[7]);
assign m2_8 = (a[2] ^ a[8]) & (b[2] ^ b[8]);
assign m2_9 = (a[2] ^ a[9]) & (b[2] ^ b[9]);
assign m2_10 = (a[2] ^ a[10]) & (b[2] ^ b[10]);
assign m2_11 = (a[2] ^ a[11]) & (b[2] ^ b[11]);
assign m2_12 = (a[2] ^ a[12]) & (b[2] ^ b[12]);
assign m2_13 = (a[2] ^ a[13]) & (b[2] ^ b[13]);
assign m2_14 = (a[2] ^ a[14]) & (b[2] ^ b[14]);
assign m2_15 = (a[2] ^ a[15]) & (b[2] ^ b[15]);
assign m2_16 = (a[2] ^ a[16]) & (b[2] ^ b[16]);
assign m2_17 = (a[2] ^ a[17]) & (b[2] ^ b[17]);
assign m2_18 = (a[2] ^ a[18]) & (b[2] ^ b[18]);
assign m2_19 = (a[2] ^ a[19]) & (b[2] ^ b[19]);
assign m2_20 = (a[2] ^ a[20]) & (b[2] ^ b[20]);
assign m2_21 = (a[2] ^ a[21]) & (b[2] ^ b[21]);
assign m2_22 = (a[2] ^ a[22]) & (b[2] ^ b[22]);
assign m2_23 = (a[2] ^ a[23]) & (b[2] ^ b[23]);
assign m2_24 = (a[2] ^ a[24]) & (b[2] ^ b[24]);
assign m2_25 = (a[2] ^ a[25]) & (b[2] ^ b[25]);
assign m3_4 = (a[3] ^ a[4]) & (b[3] ^ b[4]);
assign m3_5 = (a[3] ^ a[5]) & (b[3] ^ b[5]);
assign m3_6 = (a[3] ^ a[6]) & (b[3] ^ b[6]);
assign m3_7 = (a[3] ^ a[7]) & (b[3] ^ b[7]);
assign m3_8 = (a[3] ^ a[8]) & (b[3] ^ b[8]);
assign m3_9 = (a[3] ^ a[9]) & (b[3] ^ b[9]);
assign m3_10 = (a[3] ^ a[10]) & (b[3] ^ b[10]);
assign m3_11 = (a[3] ^ a[11]) & (b[3] ^ b[11]);
assign m3_12 = (a[3] ^ a[12]) & (b[3] ^ b[12]);
assign m3_13 = (a[3] ^ a[13]) & (b[3] ^ b[13]);
assign m3_14 = (a[3] ^ a[14]) & (b[3] ^ b[14]);
assign m3_15 = (a[3] ^ a[15]) & (b[3] ^ b[15]);
assign m3_16 = (a[3] ^ a[16]) & (b[3] ^ b[16]);
assign m3_17 = (a[3] ^ a[17]) & (b[3] ^ b[17]);
assign m3_18 = (a[3] ^ a[18]) & (b[3] ^ b[18]);
assign m3_19 = (a[3] ^ a[19]) & (b[3] ^ b[19]);
assign m3_20 = (a[3] ^ a[20]) & (b[3] ^ b[20]);
assign m3_21 = (a[3] ^ a[21]) & (b[3] ^ b[21]);
assign m3_22 = (a[3] ^ a[22]) & (b[3] ^ b[22]);
assign m3_23 = (a[3] ^ a[23]) & (b[3] ^ b[23]);
assign m3_24 = (a[3] ^ a[24]) & (b[3] ^ b[24]);
assign m3_25 = (a[3] ^ a[25]) & (b[3] ^ b[25]);
assign m4_5 = (a[4] ^ a[5]) & (b[4] ^ b[5]);
assign m4_6 = (a[4] ^ a[6]) & (b[4] ^ b[6]);
assign m4_7 = (a[4] ^ a[7]) & (b[4] ^ b[7]);
assign m4_8 = (a[4] ^ a[8]) & (b[4] ^ b[8]);
assign m4_9 = (a[4] ^ a[9]) & (b[4] ^ b[9]);
assign m4_10 = (a[4] ^ a[10]) & (b[4] ^ b[10]);
assign m4_11 = (a[4] ^ a[11]) & (b[4] ^ b[11]);
assign m4_12 = (a[4] ^ a[12]) & (b[4] ^ b[12]);
assign m4_13 = (a[4] ^ a[13]) & (b[4] ^ b[13]);
assign m4_14 = (a[4] ^ a[14]) & (b[4] ^ b[14]);
assign m4_15 = (a[4] ^ a[15]) & (b[4] ^ b[15]);
assign m4_16 = (a[4] ^ a[16]) & (b[4] ^ b[16]);
assign m4_17 = (a[4] ^ a[17]) & (b[4] ^ b[17]);
assign m4_18 = (a[4] ^ a[18]) & (b[4] ^ b[18]);
assign m4_19 = (a[4] ^ a[19]) & (b[4] ^ b[19]);
assign m4_20 = (a[4] ^ a[20]) & (b[4] ^ b[20]);
assign m4_21 = (a[4] ^ a[21]) & (b[4] ^ b[21]);
assign m4_22 = (a[4] ^ a[22]) & (b[4] ^ b[22]);
assign m4_23 = (a[4] ^ a[23]) & (b[4] ^ b[23]);
assign m4_24 = (a[4] ^ a[24]) & (b[4] ^ b[24]);
assign m4_25 = (a[4] ^ a[25]) & (b[4] ^ b[25]);
assign m5_6 = (a[5] ^ a[6]) & (b[5] ^ b[6]);
assign m5_7 = (a[5] ^ a[7]) & (b[5] ^ b[7]);
assign m5_8 = (a[5] ^ a[8]) & (b[5] ^ b[8]);
assign m5_9 = (a[5] ^ a[9]) & (b[5] ^ b[9]);
assign m5_10 = (a[5] ^ a[10]) & (b[5] ^ b[10]);
assign m5_11 = (a[5] ^ a[11]) & (b[5] ^ b[11]);
assign m5_12 = (a[5] ^ a[12]) & (b[5] ^ b[12]);
assign m5_13 = (a[5] ^ a[13]) & (b[5] ^ b[13]);
assign m5_14 = (a[5] ^ a[14]) & (b[5] ^ b[14]);
assign m5_15 = (a[5] ^ a[15]) & (b[5] ^ b[15]);
assign m5_16 = (a[5] ^ a[16]) & (b[5] ^ b[16]);
assign m5_17 = (a[5] ^ a[17]) & (b[5] ^ b[17]);
assign m5_18 = (a[5] ^ a[18]) & (b[5] ^ b[18]);
assign m5_19 = (a[5] ^ a[19]) & (b[5] ^ b[19]);
assign m5_20 = (a[5] ^ a[20]) & (b[5] ^ b[20]);
assign m5_21 = (a[5] ^ a[21]) & (b[5] ^ b[21]);
assign m5_22 = (a[5] ^ a[22]) & (b[5] ^ b[22]);
assign m5_23 = (a[5] ^ a[23]) & (b[5] ^ b[23]);
assign m5_24 = (a[5] ^ a[24]) & (b[5] ^ b[24]);
assign m5_25 = (a[5] ^ a[25]) & (b[5] ^ b[25]);
assign m6_7 = (a[6] ^ a[7]) & (b[6] ^ b[7]);
assign m6_8 = (a[6] ^ a[8]) & (b[6] ^ b[8]);
assign m6_9 = (a[6] ^ a[9]) & (b[6] ^ b[9]);
assign m6_10 = (a[6] ^ a[10]) & (b[6] ^ b[10]);
assign m6_11 = (a[6] ^ a[11]) & (b[6] ^ b[11]);
assign m6_12 = (a[6] ^ a[12]) & (b[6] ^ b[12]);
assign m6_13 = (a[6] ^ a[13]) & (b[6] ^ b[13]);
assign m6_14 = (a[6] ^ a[14]) & (b[6] ^ b[14]);
assign m6_15 = (a[6] ^ a[15]) & (b[6] ^ b[15]);
assign m6_16 = (a[6] ^ a[16]) & (b[6] ^ b[16]);
assign m6_17 = (a[6] ^ a[17]) & (b[6] ^ b[17]);
assign m6_18 = (a[6] ^ a[18]) & (b[6] ^ b[18]);
assign m6_19 = (a[6] ^ a[19]) & (b[6] ^ b[19]);
assign m6_20 = (a[6] ^ a[20]) & (b[6] ^ b[20]);
assign m6_21 = (a[6] ^ a[21]) & (b[6] ^ b[21]);
assign m6_22 = (a[6] ^ a[22]) & (b[6] ^ b[22]);
assign m6_23 = (a[6] ^ a[23]) & (b[6] ^ b[23]);
assign m6_24 = (a[6] ^ a[24]) & (b[6] ^ b[24]);
assign m6_25 = (a[6] ^ a[25]) & (b[6] ^ b[25]);
assign m7_8 = (a[7] ^ a[8]) & (b[7] ^ b[8]);
assign m7_9 = (a[7] ^ a[9]) & (b[7] ^ b[9]);
assign m7_10 = (a[7] ^ a[10]) & (b[7] ^ b[10]);
assign m7_11 = (a[7] ^ a[11]) & (b[7] ^ b[11]);
assign m7_12 = (a[7] ^ a[12]) & (b[7] ^ b[12]);
assign m7_13 = (a[7] ^ a[13]) & (b[7] ^ b[13]);
assign m7_14 = (a[7] ^ a[14]) & (b[7] ^ b[14]);
assign m7_15 = (a[7] ^ a[15]) & (b[7] ^ b[15]);
assign m7_16 = (a[7] ^ a[16]) & (b[7] ^ b[16]);
assign m7_17 = (a[7] ^ a[17]) & (b[7] ^ b[17]);
assign m7_18 = (a[7] ^ a[18]) & (b[7] ^ b[18]);
assign m7_19 = (a[7] ^ a[19]) & (b[7] ^ b[19]);
assign m7_20 = (a[7] ^ a[20]) & (b[7] ^ b[20]);
assign m7_21 = (a[7] ^ a[21]) & (b[7] ^ b[21]);
assign m7_22 = (a[7] ^ a[22]) & (b[7] ^ b[22]);
assign m7_23 = (a[7] ^ a[23]) & (b[7] ^ b[23]);
assign m7_24 = (a[7] ^ a[24]) & (b[7] ^ b[24]);
assign m7_25 = (a[7] ^ a[25]) & (b[7] ^ b[25]);
assign m8_9 = (a[8] ^ a[9]) & (b[8] ^ b[9]);
assign m8_10 = (a[8] ^ a[10]) & (b[8] ^ b[10]);
assign m8_11 = (a[8] ^ a[11]) & (b[8] ^ b[11]);
assign m8_12 = (a[8] ^ a[12]) & (b[8] ^ b[12]);
assign m8_13 = (a[8] ^ a[13]) & (b[8] ^ b[13]);
assign m8_14 = (a[8] ^ a[14]) & (b[8] ^ b[14]);
assign m8_15 = (a[8] ^ a[15]) & (b[8] ^ b[15]);
assign m8_16 = (a[8] ^ a[16]) & (b[8] ^ b[16]);
assign m8_17 = (a[8] ^ a[17]) & (b[8] ^ b[17]);
assign m8_18 = (a[8] ^ a[18]) & (b[8] ^ b[18]);
assign m8_19 = (a[8] ^ a[19]) & (b[8] ^ b[19]);
assign m8_20 = (a[8] ^ a[20]) & (b[8] ^ b[20]);
assign m8_21 = (a[8] ^ a[21]) & (b[8] ^ b[21]);
assign m8_22 = (a[8] ^ a[22]) & (b[8] ^ b[22]);
assign m8_23 = (a[8] ^ a[23]) & (b[8] ^ b[23]);
assign m8_24 = (a[8] ^ a[24]) & (b[8] ^ b[24]);
assign m8_25 = (a[8] ^ a[25]) & (b[8] ^ b[25]);
assign m9_10 = (a[9] ^ a[10]) & (b[9] ^ b[10]);
assign m9_11 = (a[9] ^ a[11]) & (b[9] ^ b[11]);
assign m9_12 = (a[9] ^ a[12]) & (b[9] ^ b[12]);
assign m9_13 = (a[9] ^ a[13]) & (b[9] ^ b[13]);
assign m9_14 = (a[9] ^ a[14]) & (b[9] ^ b[14]);
assign m9_15 = (a[9] ^ a[15]) & (b[9] ^ b[15]);
assign m9_16 = (a[9] ^ a[16]) & (b[9] ^ b[16]);
assign m9_17 = (a[9] ^ a[17]) & (b[9] ^ b[17]);
assign m9_18 = (a[9] ^ a[18]) & (b[9] ^ b[18]);
assign m9_19 = (a[9] ^ a[19]) & (b[9] ^ b[19]);
assign m9_20 = (a[9] ^ a[20]) & (b[9] ^ b[20]);
assign m9_21 = (a[9] ^ a[21]) & (b[9] ^ b[21]);
assign m9_22 = (a[9] ^ a[22]) & (b[9] ^ b[22]);
assign m9_23 = (a[9] ^ a[23]) & (b[9] ^ b[23]);
assign m9_24 = (a[9] ^ a[24]) & (b[9] ^ b[24]);
assign m9_25 = (a[9] ^ a[25]) & (b[9] ^ b[25]);
assign m10_11 = (a[10] ^ a[11]) & (b[10] ^ b[11]);
assign m10_12 = (a[10] ^ a[12]) & (b[10] ^ b[12]);
assign m10_13 = (a[10] ^ a[13]) & (b[10] ^ b[13]);
assign m10_14 = (a[10] ^ a[14]) & (b[10] ^ b[14]);
assign m10_15 = (a[10] ^ a[15]) & (b[10] ^ b[15]);
assign m10_16 = (a[10] ^ a[16]) & (b[10] ^ b[16]);
assign m10_17 = (a[10] ^ a[17]) & (b[10] ^ b[17]);
assign m10_18 = (a[10] ^ a[18]) & (b[10] ^ b[18]);
assign m10_19 = (a[10] ^ a[19]) & (b[10] ^ b[19]);
assign m10_20 = (a[10] ^ a[20]) & (b[10] ^ b[20]);
assign m10_21 = (a[10] ^ a[21]) & (b[10] ^ b[21]);
assign m10_22 = (a[10] ^ a[22]) & (b[10] ^ b[22]);
assign m10_23 = (a[10] ^ a[23]) & (b[10] ^ b[23]);
assign m10_24 = (a[10] ^ a[24]) & (b[10] ^ b[24]);
assign m10_25 = (a[10] ^ a[25]) & (b[10] ^ b[25]);
assign m11_12 = (a[11] ^ a[12]) & (b[11] ^ b[12]);
assign m11_13 = (a[11] ^ a[13]) & (b[11] ^ b[13]);
assign m11_14 = (a[11] ^ a[14]) & (b[11] ^ b[14]);
assign m11_15 = (a[11] ^ a[15]) & (b[11] ^ b[15]);
assign m11_16 = (a[11] ^ a[16]) & (b[11] ^ b[16]);
assign m11_17 = (a[11] ^ a[17]) & (b[11] ^ b[17]);
assign m11_18 = (a[11] ^ a[18]) & (b[11] ^ b[18]);
assign m11_19 = (a[11] ^ a[19]) & (b[11] ^ b[19]);
assign m11_20 = (a[11] ^ a[20]) & (b[11] ^ b[20]);
assign m11_21 = (a[11] ^ a[21]) & (b[11] ^ b[21]);
assign m11_22 = (a[11] ^ a[22]) & (b[11] ^ b[22]);
assign m11_23 = (a[11] ^ a[23]) & (b[11] ^ b[23]);
assign m11_24 = (a[11] ^ a[24]) & (b[11] ^ b[24]);
assign m11_25 = (a[11] ^ a[25]) & (b[11] ^ b[25]);
assign m12_13 = (a[12] ^ a[13]) & (b[12] ^ b[13]);
assign m12_14 = (a[12] ^ a[14]) & (b[12] ^ b[14]);
assign m12_15 = (a[12] ^ a[15]) & (b[12] ^ b[15]);
assign m12_16 = (a[12] ^ a[16]) & (b[12] ^ b[16]);
assign m12_17 = (a[12] ^ a[17]) & (b[12] ^ b[17]);
assign m12_18 = (a[12] ^ a[18]) & (b[12] ^ b[18]);
assign m12_19 = (a[12] ^ a[19]) & (b[12] ^ b[19]);
assign m12_20 = (a[12] ^ a[20]) & (b[12] ^ b[20]);
assign m12_21 = (a[12] ^ a[21]) & (b[12] ^ b[21]);
assign m12_22 = (a[12] ^ a[22]) & (b[12] ^ b[22]);
assign m12_23 = (a[12] ^ a[23]) & (b[12] ^ b[23]);
assign m12_24 = (a[12] ^ a[24]) & (b[12] ^ b[24]);
assign m12_25 = (a[12] ^ a[25]) & (b[12] ^ b[25]);
assign m13_14 = (a[13] ^ a[14]) & (b[13] ^ b[14]);
assign m13_15 = (a[13] ^ a[15]) & (b[13] ^ b[15]);
assign m13_16 = (a[13] ^ a[16]) & (b[13] ^ b[16]);
assign m13_17 = (a[13] ^ a[17]) & (b[13] ^ b[17]);
assign m13_18 = (a[13] ^ a[18]) & (b[13] ^ b[18]);
assign m13_19 = (a[13] ^ a[19]) & (b[13] ^ b[19]);
assign m13_20 = (a[13] ^ a[20]) & (b[13] ^ b[20]);
assign m13_21 = (a[13] ^ a[21]) & (b[13] ^ b[21]);
assign m13_22 = (a[13] ^ a[22]) & (b[13] ^ b[22]);
assign m13_23 = (a[13] ^ a[23]) & (b[13] ^ b[23]);
assign m13_24 = (a[13] ^ a[24]) & (b[13] ^ b[24]);
assign m13_25 = (a[13] ^ a[25]) & (b[13] ^ b[25]);
assign m14_15 = (a[14] ^ a[15]) & (b[14] ^ b[15]);
assign m14_16 = (a[14] ^ a[16]) & (b[14] ^ b[16]);
assign m14_17 = (a[14] ^ a[17]) & (b[14] ^ b[17]);
assign m14_18 = (a[14] ^ a[18]) & (b[14] ^ b[18]);
assign m14_19 = (a[14] ^ a[19]) & (b[14] ^ b[19]);
assign m14_20 = (a[14] ^ a[20]) & (b[14] ^ b[20]);
assign m14_21 = (a[14] ^ a[21]) & (b[14] ^ b[21]);
assign m14_22 = (a[14] ^ a[22]) & (b[14] ^ b[22]);
assign m14_23 = (a[14] ^ a[23]) & (b[14] ^ b[23]);
assign m14_24 = (a[14] ^ a[24]) & (b[14] ^ b[24]);
assign m14_25 = (a[14] ^ a[25]) & (b[14] ^ b[25]);
assign m15_16 = (a[15] ^ a[16]) & (b[15] ^ b[16]);
assign m15_17 = (a[15] ^ a[17]) & (b[15] ^ b[17]);
assign m15_18 = (a[15] ^ a[18]) & (b[15] ^ b[18]);
assign m15_19 = (a[15] ^ a[19]) & (b[15] ^ b[19]);
assign m15_20 = (a[15] ^ a[20]) & (b[15] ^ b[20]);
assign m15_21 = (a[15] ^ a[21]) & (b[15] ^ b[21]);
assign m15_22 = (a[15] ^ a[22]) & (b[15] ^ b[22]);
assign m15_23 = (a[15] ^ a[23]) & (b[15] ^ b[23]);
assign m15_24 = (a[15] ^ a[24]) & (b[15] ^ b[24]);
assign m15_25 = (a[15] ^ a[25]) & (b[15] ^ b[25]);
assign m16_17 = (a[16] ^ a[17]) & (b[16] ^ b[17]);
assign m16_18 = (a[16] ^ a[18]) & (b[16] ^ b[18]);
assign m16_19 = (a[16] ^ a[19]) & (b[16] ^ b[19]);
assign m16_20 = (a[16] ^ a[20]) & (b[16] ^ b[20]);
assign m16_21 = (a[16] ^ a[21]) & (b[16] ^ b[21]);
assign m16_22 = (a[16] ^ a[22]) & (b[16] ^ b[22]);
assign m16_23 = (a[16] ^ a[23]) & (b[16] ^ b[23]);
assign m16_24 = (a[16] ^ a[24]) & (b[16] ^ b[24]);
assign m16_25 = (a[16] ^ a[25]) & (b[16] ^ b[25]);
assign m17_18 = (a[17] ^ a[18]) & (b[17] ^ b[18]);
assign m17_19 = (a[17] ^ a[19]) & (b[17] ^ b[19]);
assign m17_20 = (a[17] ^ a[20]) & (b[17] ^ b[20]);
assign m17_21 = (a[17] ^ a[21]) & (b[17] ^ b[21]);
assign m17_22 = (a[17] ^ a[22]) & (b[17] ^ b[22]);
assign m17_23 = (a[17] ^ a[23]) & (b[17] ^ b[23]);
assign m17_24 = (a[17] ^ a[24]) & (b[17] ^ b[24]);
assign m17_25 = (a[17] ^ a[25]) & (b[17] ^ b[25]);
assign m18_19 = (a[18] ^ a[19]) & (b[18] ^ b[19]);
assign m18_20 = (a[18] ^ a[20]) & (b[18] ^ b[20]);
assign m18_21 = (a[18] ^ a[21]) & (b[18] ^ b[21]);
assign m18_22 = (a[18] ^ a[22]) & (b[18] ^ b[22]);
assign m18_23 = (a[18] ^ a[23]) & (b[18] ^ b[23]);
assign m18_24 = (a[18] ^ a[24]) & (b[18] ^ b[24]);
assign m18_25 = (a[18] ^ a[25]) & (b[18] ^ b[25]);
assign m19_20 = (a[19] ^ a[20]) & (b[19] ^ b[20]);
assign m19_21 = (a[19] ^ a[21]) & (b[19] ^ b[21]);
assign m19_22 = (a[19] ^ a[22]) & (b[19] ^ b[22]);
assign m19_23 = (a[19] ^ a[23]) & (b[19] ^ b[23]);
assign m19_24 = (a[19] ^ a[24]) & (b[19] ^ b[24]);
assign m19_25 = (a[19] ^ a[25]) & (b[19] ^ b[25]);
assign m20_21 = (a[20] ^ a[21]) & (b[20] ^ b[21]);
assign m20_22 = (a[20] ^ a[22]) & (b[20] ^ b[22]);
assign m20_23 = (a[20] ^ a[23]) & (b[20] ^ b[23]);
assign m20_24 = (a[20] ^ a[24]) & (b[20] ^ b[24]);
assign m20_25 = (a[20] ^ a[25]) & (b[20] ^ b[25]);
assign m21_22 = (a[21] ^ a[22]) & (b[21] ^ b[22]);
assign m21_23 = (a[21] ^ a[23]) & (b[21] ^ b[23]);
assign m21_24 = (a[21] ^ a[24]) & (b[21] ^ b[24]);
assign m21_25 = (a[21] ^ a[25]) & (b[21] ^ b[25]);
assign m22_23 = (a[22] ^ a[23]) & (b[22] ^ b[23]);
assign m22_24 = (a[22] ^ a[24]) & (b[22] ^ b[24]);
assign m22_25 = (a[22] ^ a[25]) & (b[22] ^ b[25]);
assign m23_24 = (a[23] ^ a[24]) & (b[23] ^ b[24]);
assign m23_25 = (a[23] ^ a[25]) & (b[23] ^ b[25]);
assign m24_25 = (a[24] ^ a[25]) & (b[24] ^ b[25]);
assign d[0] = m0;
assign d[1] = m0_1 ^ m0 ^ m1;
assign d[2] = m0_2 ^ m0 ^ m1 ^ m2;
assign d[3] = m0_3 ^ m1_2 ^ m0 ^ m1 ^ m2 ^ m3;
assign d[4] = m0_4 ^ m1_3 ^ m0 ^ m1 ^ m2 ^ m3 ^ m4;
assign d[5] = m0_5 ^ m1_4 ^ m2_3 ^ m0 ^ m1 ^ m2 ^ m3 ^ m4 ^ m5;
assign d[6] = m0_6 ^ m1_5 ^ m2_4 ^ m0 ^ m1 ^ m2 ^ m3 ^ m4 ^ m5 ^ m6;
assign d[7] = m0_7 ^ m1_6 ^ m2_5 ^ m3_4 ^ m0 ^ m1 ^ m2 ^ m3 ^ m4 ^ m5 ^ m6 ^ m7;
assign d[8] = m0_8 ^ m1_7 ^ m2_6 ^ m3_5 ^ m0 ^ m1 ^ m2 ^ m3 ^ m4 ^ m5 ^ m6 ^ m7 ^ m8;
assign d[9] = m0_9 ^ m1_8 ^ m2_7 ^ m3_6 ^ m4_5 ^ m0 ^ m1 ^ m2 ^ m3 ^ m4 ^ m5 ^ m6 ^ m7 ^ m8 ^ m9;
assign d[10] = m0_10 ^ m1_9 ^ m2_8 ^ m3_7 ^ m4_6 ^ m0 ^ m1 ^ m2 ^ m3 ^ m4 ^ m5 ^ m6 ^ m7 ^ m8 ^ m9 ^ m10;
assign d[11] = m0_11 ^ m1_10 ^ m2_9 ^ m3_8 ^ m4_7 ^ m5_6 ^ m0 ^ m1 ^ m2 ^ m3 ^ m4 ^ m5 ^ m6 ^ m7 ^ m8 ^ m9 ^ m10 ^ m11;
assign d[12] = m0_12 ^ m1_11 ^ m2_10 ^ m3_9 ^ m4_8 ^ m5_7 ^ m0 ^ m1 ^ m2 ^ m3 ^ m4 ^ m5 ^ m6 ^ m7 ^ m8 ^ m9 ^ m10 ^ m11 ^ m12;
assign d[13] = m0_13 ^ m1_12 ^ m2_11 ^ m3_10 ^ m4_9 ^ m5_8 ^ m6_7 ^ m0 ^ m1 ^ m2 ^ m3 ^ m4 ^ m5 ^ m6 ^ m7 ^ m8 ^ m9 ^ m10 ^ m11 ^ m12 ^ m13;
assign d[14] = m0_14 ^ m1_13 ^ m2_12 ^ m3_11 ^ m4_10 ^ m5_9 ^ m6_8 ^ m0 ^ m1 ^ m2 ^ m3 ^ m4 ^ m5 ^ m6 ^ m7 ^ m8 ^ m9 ^ m10 ^ m11 ^ m12 ^ m13 ^ m14;
assign d[15] = m0_15 ^ m1_14 ^ m2_13 ^ m3_12 ^ m4_11 ^ m5_10 ^ m6_9 ^ m7_8 ^ m0 ^ m1 ^ m2 ^ m3 ^ m4 ^ m5 ^ m6 ^ m7 ^ m8 ^ m9 ^ m10 ^ m11 ^ m12 ^ m13 ^ m14 ^ m15;
assign d[16] = m0_16 ^ m1_15 ^ m2_14 ^ m3_13 ^ m4_12 ^ m5_11 ^ m6_10 ^ m7_9 ^ m0 ^ m1 ^ m2 ^ m3 ^ m4 ^ m5 ^ m6 ^ m7 ^ m8 ^ m9 ^ m10 ^ m11 ^ m12 ^ m13 ^ m14 ^ m15 ^ m16;
assign d[17] = m0_17 ^ m1_16 ^ m2_15 ^ m3_14 ^ m4_13 ^ m5_12 ^ m6_11 ^ m7_10 ^ m8_9 ^ m0 ^ m1 ^ m2 ^ m3 ^ m4 ^ m5 ^ m6 ^ m7 ^ m8 ^ m9 ^ m10 ^ m11 ^ m12 ^ m13 ^ m14 ^ m15 ^ m16 ^ m17;
assign d[18] = m0_18 ^ m1_17 ^ m2_16 ^ m3_15 ^ m4_14 ^ m5_13 ^ m6_12 ^ m7_11 ^ m8_10 ^ m0 ^ m1 ^ m2 ^ m3 ^ m4 ^ m5 ^ m6 ^ m7 ^ m8 ^ m9 ^ m10 ^ m11 ^ m12 ^ m13 ^ m14 ^ m15 ^ m16 ^ m17 ^ m18;
assign d[19] = m0_19 ^ m1_18 ^ m2_17 ^ m3_16 ^ m4_15 ^ m5_14 ^ m6_13 ^ m7_12 ^ m8_11 ^ m9_10 ^ m0 ^ m1 ^ m2 ^ m3 ^ m4 ^ m5 ^ m6 ^ m7 ^ m8 ^ m9 ^ m10 ^ m11 ^ m12 ^ m13 ^ m14 ^ m15 ^ m16 ^ m17 ^ m18 ^ m19;
assign d[20] = m0_20 ^ m1_19 ^ m2_18 ^ m3_17 ^ m4_16 ^ m5_15 ^ m6_14 ^ m7_13 ^ m8_12 ^ m9_11 ^ m0 ^ m1 ^ m2 ^ m3 ^ m4 ^ m5 ^ m6 ^ m7 ^ m8 ^ m9 ^ m10 ^ m11 ^ m12 ^ m13 ^ m14 ^ m15 ^ m16 ^ m17 ^ m18 ^ m19 ^ m20;
assign d[21] = m0_21 ^ m1_20 ^ m2_19 ^ m3_18 ^ m4_17 ^ m5_16 ^ m6_15 ^ m7_14 ^ m8_13 ^ m9_12 ^ m10_11 ^ m0 ^ m1 ^ m2 ^ m3 ^ m4 ^ m5 ^ m6 ^ m7 ^ m8 ^ m9 ^ m10 ^ m11 ^ m12 ^ m13 ^ m14 ^ m15 ^ m16 ^ m17 ^ m18 ^ m19 ^ m20 ^ m21;
assign d[22] = m0_22 ^ m1_21 ^ m2_20 ^ m3_19 ^ m4_18 ^ m5_17 ^ m6_16 ^ m7_15 ^ m8_14 ^ m9_13 ^ m10_12 ^ m0 ^ m1 ^ m2 ^ m3 ^ m4 ^ m5 ^ m6 ^ m7 ^ m8 ^ m9 ^ m10 ^ m11 ^ m12 ^ m13 ^ m14 ^ m15 ^ m16 ^ m17 ^ m18 ^ m19 ^ m20 ^ m21 ^ m22;
assign d[23] = m0_23 ^ m1_22 ^ m2_21 ^ m3_20 ^ m4_19 ^ m5_18 ^ m6_17 ^ m7_16 ^ m8_15 ^ m9_14 ^ m10_13 ^ m11_12 ^ m0 ^ m1 ^ m2 ^ m3 ^ m4 ^ m5 ^ m6 ^ m7 ^ m8 ^ m9 ^ m10 ^ m11 ^ m12 ^ m13 ^ m14 ^ m15 ^ m16 ^ m17 ^ m18 ^ m19 ^ m20 ^ m21 ^ m22 ^ m23;
assign d[24] = m0_24 ^ m1_23 ^ m2_22 ^ m3_21 ^ m4_20 ^ m5_19 ^ m6_18 ^ m7_17 ^ m8_16 ^ m9_15 ^ m10_14 ^ m11_13 ^ m0 ^ m1 ^ m2 ^ m3 ^ m4 ^ m5 ^ m6 ^ m7 ^ m8 ^ m9 ^ m10 ^ m11 ^ m12 ^ m13 ^ m14 ^ m15 ^ m16 ^ m17 ^ m18 ^ m19 ^ m20 ^ m21 ^ m22 ^ m23 ^ m24;
assign d[25] = m0_25 ^ m1_24 ^ m2_23 ^ m3_22 ^ m4_21 ^ m5_20 ^ m6_19 ^ m7_18 ^ m8_17 ^ m9_16 ^ m10_15 ^ m11_14 ^ m12_13 ^ m0 ^ m1 ^ m2 ^ m3 ^ m4 ^ m5 ^ m6 ^ m7 ^ m8 ^ m9 ^ m10 ^ m11 ^ m12 ^ m13 ^ m14 ^ m15 ^ m16 ^ m17 ^ m18 ^ m19 ^ m20 ^ m21 ^ m22 ^ m23 ^ m24 ^ m25;
assign d[26] = m1_25 ^ m2_24 ^ m3_23 ^ m4_22 ^ m5_21 ^ m6_20 ^ m7_19 ^ m8_18 ^ m9_17 ^ m10_16 ^ m11_15 ^ m12_14 ^ m1 ^ m2 ^ m3 ^ m4 ^ m5 ^ m6 ^ m7 ^ m8 ^ m9 ^ m10 ^ m11 ^ m12 ^ m13 ^ m14 ^ m15 ^ m16 ^ m17 ^ m18 ^ m19 ^ m20 ^ m21 ^ m22 ^ m23 ^ m24 ^ m25;
assign d[27] = m2_25 ^ m3_24 ^ m4_23 ^ m5_22 ^ m6_21 ^ m7_20 ^ m8_19 ^ m9_18 ^ m10_17 ^ m11_16 ^ m12_15 ^ m13_14 ^ m2 ^ m3 ^ m4 ^ m5 ^ m6 ^ m7 ^ m8 ^ m9 ^ m10 ^ m11 ^ m12 ^ m13 ^ m14 ^ m15 ^ m16 ^ m17 ^ m18 ^ m19 ^ m20 ^ m21 ^ m22 ^ m23 ^ m24 ^ m25;
assign d[28] = m3_25 ^ m4_24 ^ m5_23 ^ m6_22 ^ m7_21 ^ m8_20 ^ m9_19 ^ m10_18 ^ m11_17 ^ m12_16 ^ m13_15 ^ m3 ^ m4 ^ m5 ^ m6 ^ m7 ^ m8 ^ m9 ^ m10 ^ m11 ^ m12 ^ m13 ^ m14 ^ m15 ^ m16 ^ m17 ^ m18 ^ m19 ^ m20 ^ m21 ^ m22 ^ m23 ^ m24 ^ m25;
assign d[29] = m4_25 ^ m5_24 ^ m6_23 ^ m7_22 ^ m8_21 ^ m9_20 ^ m10_19 ^ m11_18 ^ m12_17 ^ m13_16 ^ m14_15 ^ m4 ^ m5 ^ m6 ^ m7 ^ m8 ^ m9 ^ m10 ^ m11 ^ m12 ^ m13 ^ m14 ^ m15 ^ m16 ^ m17 ^ m18 ^ m19 ^ m20 ^ m21 ^ m22 ^ m23 ^ m24 ^ m25;
assign d[30] = m5_25 ^ m6_24 ^ m7_23 ^ m8_22 ^ m9_21 ^ m10_20 ^ m11_19 ^ m12_18 ^ m13_17 ^ m14_16 ^ m5 ^ m6 ^ m7 ^ m8 ^ m9 ^ m10 ^ m11 ^ m12 ^ m13 ^ m14 ^ m15 ^ m16 ^ m17 ^ m18 ^ m19 ^ m20 ^ m21 ^ m22 ^ m23 ^ m24 ^ m25;
assign d[31] = m6_25 ^ m7_24 ^ m8_23 ^ m9_22 ^ m10_21 ^ m11_20 ^ m12_19 ^ m13_18 ^ m14_17 ^ m15_16 ^ m6 ^ m7 ^ m8 ^ m9 ^ m10 ^ m11 ^ m12 ^ m13 ^ m14 ^ m15 ^ m16 ^ m17 ^ m18 ^ m19 ^ m20 ^ m21 ^ m22 ^ m23 ^ m24 ^ m25;
assign d[32] = m7_25 ^ m8_24 ^ m9_23 ^ m10_22 ^ m11_21 ^ m12_20 ^ m13_19 ^ m14_18 ^ m15_17 ^ m7 ^ m8 ^ m9 ^ m10 ^ m11 ^ m12 ^ m13 ^ m14 ^ m15 ^ m16 ^ m17 ^ m18 ^ m19 ^ m20 ^ m21 ^ m22 ^ m23 ^ m24 ^ m25;
assign d[33] = m8_25 ^ m9_24 ^ m10_23 ^ m11_22 ^ m12_21 ^ m13_20 ^ m14_19 ^ m15_18 ^ m16_17 ^ m8 ^ m9 ^ m10 ^ m11 ^ m12 ^ m13 ^ m14 ^ m15 ^ m16 ^ m17 ^ m18 ^ m19 ^ m20 ^ m21 ^ m22 ^ m23 ^ m24 ^ m25;
assign d[34] = m9_25 ^ m10_24 ^ m11_23 ^ m12_22 ^ m13_21 ^ m14_20 ^ m15_19 ^ m16_18 ^ m9 ^ m10 ^ m11 ^ m12 ^ m13 ^ m14 ^ m15 ^ m16 ^ m17 ^ m18 ^ m19 ^ m20 ^ m21 ^ m22 ^ m23 ^ m24 ^ m25;
assign d[35] = m10_25 ^ m11_24 ^ m12_23 ^ m13_22 ^ m14_21 ^ m15_20 ^ m16_19 ^ m17_18 ^ m10 ^ m11 ^ m12 ^ m13 ^ m14 ^ m15 ^ m16 ^ m17 ^ m18 ^ m19 ^ m20 ^ m21 ^ m22 ^ m23 ^ m24 ^ m25;
assign d[36] = m11_25 ^ m12_24 ^ m13_23 ^ m14_22 ^ m15_21 ^ m16_20 ^ m17_19 ^ m11 ^ m12 ^ m13 ^ m14 ^ m15 ^ m16 ^ m17 ^ m18 ^ m19 ^ m20 ^ m21 ^ m22 ^ m23 ^ m24 ^ m25;
assign d[37] = m12_25 ^ m13_24 ^ m14_23 ^ m15_22 ^ m16_21 ^ m17_20 ^ m18_19 ^ m12 ^ m13 ^ m14 ^ m15 ^ m16 ^ m17 ^ m18 ^ m19 ^ m20 ^ m21 ^ m22 ^ m23 ^ m24 ^ m25;
assign d[38] = m13_25 ^ m14_24 ^ m15_23 ^ m16_22 ^ m17_21 ^ m18_20 ^ m13 ^ m14 ^ m15 ^ m16 ^ m17 ^ m18 ^ m19 ^ m20 ^ m21 ^ m22 ^ m23 ^ m24 ^ m25;
assign d[39] = m14_25 ^ m15_24 ^ m16_23 ^ m17_22 ^ m18_21 ^ m19_20 ^ m14 ^ m15 ^ m16 ^ m17 ^ m18 ^ m19 ^ m20 ^ m21 ^ m22 ^ m23 ^ m24 ^ m25;
assign d[40] = m15_25 ^ m16_24 ^ m17_23 ^ m18_22 ^ m19_21 ^ m15 ^ m16 ^ m17 ^ m18 ^ m19 ^ m20 ^ m21 ^ m22 ^ m23 ^ m24 ^ m25;
assign d[41] = m16_25 ^ m17_24 ^ m18_23 ^ m19_22 ^ m20_21 ^ m16 ^ m17 ^ m18 ^ m19 ^ m20 ^ m21 ^ m22 ^ m23 ^ m24 ^ m25;
assign d[42] = m17_25 ^ m18_24 ^ m19_23 ^ m20_22 ^ m17 ^ m18 ^ m19 ^ m20 ^ m21 ^ m22 ^ m23 ^ m24 ^ m25;
assign d[43] = m18_25 ^ m19_24 ^ m20_23 ^ m21_22 ^ m18 ^ m19 ^ m20 ^ m21 ^ m22 ^ m23 ^ m24 ^ m25;
assign d[44] = m19_25 ^ m20_24 ^ m21_23 ^ m19 ^ m20 ^ m21 ^ m22 ^ m23 ^ m24 ^ m25;
assign d[45] = m20_25 ^ m21_24 ^ m22_23 ^ m20 ^ m21 ^ m22 ^ m23 ^ m24 ^ m25;
assign d[46] = m21_25 ^ m22_24 ^ m21 ^ m22 ^ m23 ^ m24 ^ m25;
assign d[47] = m22_25 ^ m23_24 ^ m22 ^ m23 ^ m24 ^ m25;
assign d[48] = m23_25 ^ m23 ^ m24 ^ m25;
assign d[49] = m24_25 ^ m24 ^ m25;
assign d[50] = m25;
endmodule
`endif
