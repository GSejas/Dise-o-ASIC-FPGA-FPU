`ifndef __POW_2P1__
`define __POW_2P1__
module squarer(a, d);

input wire [232:0] a;
output wire [232:0] d;

assign d[0] = a[0] ^ a[196];
assign d[1] = a[117];
assign d[2] = a[1] ^ a[197];
assign d[3] = a[118];
assign d[4] = a[2] ^ a[198];
assign d[5] = a[119];
assign d[6] = a[3] ^ a[199];
assign d[7] = a[120];
assign d[8] = a[4] ^ a[200];
assign d[9] = a[121];
assign d[10] = a[5] ^ a[201];
assign d[11] = a[122];
assign d[12] = a[6] ^ a[202];
assign d[13] = a[123];
assign d[14] = a[7] ^ a[203];
assign d[15] = a[124];
assign d[16] = a[8] ^ a[204];
assign d[17] = a[125];
assign d[18] = a[9] ^ a[205];
assign d[19] = a[126];
assign d[20] = a[10] ^ a[206];
assign d[21] = a[127];
assign d[22] = a[11] ^ a[207];
assign d[23] = a[128];
assign d[24] = a[12] ^ a[208];
assign d[25] = a[129];
assign d[26] = a[13] ^ a[209];
assign d[27] = a[130];
assign d[28] = a[14] ^ a[210];
assign d[29] = a[131];
assign d[30] = a[15] ^ a[211];
assign d[31] = a[132];
assign d[32] = a[16] ^ a[212];
assign d[33] = a[133];
assign d[34] = a[17] ^ a[213];
assign d[35] = a[134];
assign d[36] = a[18] ^ a[214];
assign d[37] = a[135];
assign d[38] = a[19] ^ a[215];
assign d[39] = a[136];
assign d[40] = a[20] ^ a[216];
assign d[41] = a[137];
assign d[42] = a[21] ^ a[217];
assign d[43] = a[138];
assign d[44] = a[22] ^ a[218];
assign d[45] = a[139];
assign d[46] = a[23] ^ a[219];
assign d[47] = a[140];
assign d[48] = a[24] ^ a[220];
assign d[49] = a[141];
assign d[50] = a[25] ^ a[221];
assign d[51] = a[142];
assign d[52] = a[26] ^ a[222];
assign d[53] = a[143];
assign d[54] = a[27] ^ a[223];
assign d[55] = a[144];
assign d[56] = a[28] ^ a[224];
assign d[57] = a[145];
assign d[58] = a[29] ^ a[225];
assign d[59] = a[146];
assign d[60] = a[30] ^ a[226];
assign d[61] = a[147];
assign d[62] = a[31] ^ a[227];
assign d[63] = a[148];
assign d[64] = a[32] ^ a[228];
assign d[65] = a[149];
assign d[66] = a[33] ^ a[229];
assign d[67] = a[150];
assign d[68] = a[34] ^ a[230];
assign d[69] = a[151];
assign d[70] = a[35] ^ a[231];
assign d[71] = a[152];
assign d[72] = a[36] ^ a[232];
assign d[73] = a[153];
assign d[74] = a[37] ^ a[196];
assign d[75] = a[117] ^ a[154];
assign d[76] = a[38] ^ a[197];
assign d[77] = a[118] ^ a[155];
assign d[78] = a[39] ^ a[198];
assign d[79] = a[119] ^ a[156];
assign d[80] = a[40] ^ a[199];
assign d[81] = a[120] ^ a[157];
assign d[82] = a[41] ^ a[200];
assign d[83] = a[121] ^ a[158];
assign d[84] = a[42] ^ a[201];
assign d[85] = a[122] ^ a[159];
assign d[86] = a[43] ^ a[202];
assign d[87] = a[123] ^ a[160];
assign d[88] = a[44] ^ a[203];
assign d[89] = a[124] ^ a[161];
assign d[90] = a[45] ^ a[204];
assign d[91] = a[125] ^ a[162];
assign d[92] = a[46] ^ a[205];
assign d[93] = a[126] ^ a[163];
assign d[94] = a[47] ^ a[206];
assign d[95] = a[127] ^ a[164];
assign d[96] = a[48] ^ a[207];
assign d[97] = a[128] ^ a[165];
assign d[98] = a[49] ^ a[208];
assign d[99] = a[129] ^ a[166];
assign d[100] = a[50] ^ a[209];
assign d[101] = a[130] ^ a[167];
assign d[102] = a[51] ^ a[210];
assign d[103] = a[131] ^ a[168];
assign d[104] = a[52] ^ a[211];
assign d[105] = a[132] ^ a[169];
assign d[106] = a[53] ^ a[212];
assign d[107] = a[133] ^ a[170];
assign d[108] = a[54] ^ a[213];
assign d[109] = a[134] ^ a[171];
assign d[110] = a[55] ^ a[214];
assign d[111] = a[135] ^ a[172];
assign d[112] = a[56] ^ a[215];
assign d[113] = a[136] ^ a[173];
assign d[114] = a[57] ^ a[216];
assign d[115] = a[137] ^ a[174];
assign d[116] = a[58] ^ a[217];
assign d[117] = a[138] ^ a[175];
assign d[118] = a[59] ^ a[218];
assign d[119] = a[139] ^ a[176];
assign d[120] = a[60] ^ a[219];
assign d[121] = a[140] ^ a[177];
assign d[122] = a[61] ^ a[220];
assign d[123] = a[141] ^ a[178];
assign d[124] = a[62] ^ a[221];
assign d[125] = a[142] ^ a[179];
assign d[126] = a[63] ^ a[222];
assign d[127] = a[143] ^ a[180];
assign d[128] = a[64] ^ a[223];
assign d[129] = a[144] ^ a[181];
assign d[130] = a[65] ^ a[224];
assign d[131] = a[145] ^ a[182];
assign d[132] = a[66] ^ a[225];
assign d[133] = a[146] ^ a[183];
assign d[134] = a[67] ^ a[226];
assign d[135] = a[147] ^ a[184];
assign d[136] = a[68] ^ a[227];
assign d[137] = a[148] ^ a[185];
assign d[138] = a[69] ^ a[228];
assign d[139] = a[149] ^ a[186];
assign d[140] = a[70] ^ a[229];
assign d[141] = a[150] ^ a[187];
assign d[142] = a[71] ^ a[230];
assign d[143] = a[151] ^ a[188];
assign d[144] = a[72] ^ a[231];
assign d[145] = a[152] ^ a[189];
assign d[146] = a[73] ^ a[232];
assign d[147] = a[153] ^ a[190];
assign d[148] = a[74];
assign d[149] = a[154] ^ a[191];
assign d[150] = a[75];
assign d[151] = a[155] ^ a[192];
assign d[152] = a[76];
assign d[153] = a[156] ^ a[193];
assign d[154] = a[77];
assign d[155] = a[157] ^ a[194];
assign d[156] = a[78];
assign d[157] = a[158] ^ a[195];
assign d[158] = a[79];
assign d[159] = a[159] ^ a[196];
assign d[160] = a[80];
assign d[161] = a[160] ^ a[197];
assign d[162] = a[81];
assign d[163] = a[161] ^ a[198];
assign d[164] = a[82];
assign d[165] = a[162] ^ a[199];
assign d[166] = a[83];
assign d[167] = a[163] ^ a[200];
assign d[168] = a[84];
assign d[169] = a[164] ^ a[201];
assign d[170] = a[85];
assign d[171] = a[165] ^ a[202];
assign d[172] = a[86];
assign d[173] = a[166] ^ a[203];
assign d[174] = a[87];
assign d[175] = a[167] ^ a[204];
assign d[176] = a[88];
assign d[177] = a[168] ^ a[205];
assign d[178] = a[89];
assign d[179] = a[169] ^ a[206];
assign d[180] = a[90];
assign d[181] = a[170] ^ a[207];
assign d[182] = a[91];
assign d[183] = a[171] ^ a[208];
assign d[184] = a[92];
assign d[185] = a[172] ^ a[209];
assign d[186] = a[93];
assign d[187] = a[173] ^ a[210];
assign d[188] = a[94];
assign d[189] = a[174] ^ a[211];
assign d[190] = a[95];
assign d[191] = a[175] ^ a[212];
assign d[192] = a[96];
assign d[193] = a[176] ^ a[213];
assign d[194] = a[97];
assign d[195] = a[177] ^ a[214];
assign d[196] = a[98];
assign d[197] = a[178] ^ a[215];
assign d[198] = a[99];
assign d[199] = a[179] ^ a[216];
assign d[200] = a[100];
assign d[201] = a[180] ^ a[217];
assign d[202] = a[101];
assign d[203] = a[181] ^ a[218];
assign d[204] = a[102];
assign d[205] = a[182] ^ a[219];
assign d[206] = a[103];
assign d[207] = a[183] ^ a[220];
assign d[208] = a[104];
assign d[209] = a[184] ^ a[221];
assign d[210] = a[105];
assign d[211] = a[185] ^ a[222];
assign d[212] = a[106];
assign d[213] = a[186] ^ a[223];
assign d[214] = a[107];
assign d[215] = a[187] ^ a[224];
assign d[216] = a[108];
assign d[217] = a[188] ^ a[225];
assign d[218] = a[109];
assign d[219] = a[189] ^ a[226];
assign d[220] = a[110];
assign d[221] = a[190] ^ a[227];
assign d[222] = a[111];
assign d[223] = a[191] ^ a[228];
assign d[224] = a[112];
assign d[225] = a[192] ^ a[229];
assign d[226] = a[113];
assign d[227] = a[193] ^ a[230];
assign d[228] = a[114];
assign d[229] = a[194] ^ a[231];
assign d[230] = a[115];
assign d[231] = a[195] ^ a[232];
assign d[232] = a[116];
endmodule
`endif
